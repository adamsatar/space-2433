`timescale 1ns / 1ps

module alien_rom(
input [9:0] address,
output reg [7:0] rgb_data
    );
(* rom_style = "block" *)


always @*
case(address)
10'd0   : rgb_data = 0;
10'd1   : rgb_data = 0;
10'd2   : rgb_data = 0;
10'd3   : rgb_data = 0;
10'd4   : rgb_data = 0;
10'd5   : rgb_data = 0;
10'd6   : rgb_data = 0;
10'd7   : rgb_data = 0;
10'd8   : rgb_data = 0;
10'd9   : rgb_data = 0;
10'd10  : rgb_data = 0;
10'd11  : rgb_data = 0;
10'd12  : rgb_data = 236;
10'd13  : rgb_data = 236;
10'd14  : rgb_data = 236;
10'd15  : rgb_data = 236;
10'd16  : rgb_data = 236;
10'd17  : rgb_data = 236;
10'd18  : rgb_data = 236;
10'd19  : rgb_data = 236;
10'd20  : rgb_data = 0;
10'd21  : rgb_data = 0;
10'd22  : rgb_data = 0;
10'd23  : rgb_data = 0;
10'd24  : rgb_data = 0;
10'd25  : rgb_data = 0;
10'd26  : rgb_data = 0;
10'd27  : rgb_data = 0;
10'd28  : rgb_data = 0;
10'd29  : rgb_data = 0;
10'd30  : rgb_data = 0;
10'd31  : rgb_data = 0;
10'd32  : rgb_data = 0;
10'd33  : rgb_data = 0;
10'd34  : rgb_data = 0;
10'd35  : rgb_data = 0;
10'd36  : rgb_data = 0;
10'd37  : rgb_data = 0;
10'd38  : rgb_data = 0;
10'd39  : rgb_data = 0;
10'd40  : rgb_data = 0;
10'd41  : rgb_data = 0;
10'd42  : rgb_data = 0;
10'd43  : rgb_data = 0;
10'd44  : rgb_data = 236;
10'd45  : rgb_data = 236;
10'd46  : rgb_data = 236;
10'd47  : rgb_data = 236;
10'd48  : rgb_data = 236;
10'd49  : rgb_data = 236;
10'd50  : rgb_data = 236;
10'd51  : rgb_data = 236;
10'd52  : rgb_data = 0;
10'd53  : rgb_data = 0;
10'd54  : rgb_data = 0;
10'd55  : rgb_data = 0;
10'd56  : rgb_data = 0;
10'd57  : rgb_data = 0;
10'd58  : rgb_data = 0;
10'd59  : rgb_data = 0;
10'd60  : rgb_data = 0;
10'd61  : rgb_data = 0;
10'd62  : rgb_data = 0;
10'd63  : rgb_data = 0;
10'd64  : rgb_data = 0;
10'd65  : rgb_data = 0;
10'd66  : rgb_data = 0;
10'd67  : rgb_data = 0;
10'd68  : rgb_data = 0;
10'd69  : rgb_data = 0;
10'd70  : rgb_data = 0;
10'd71  : rgb_data = 0;
10'd72  : rgb_data = 0;
10'd73  : rgb_data = 0;
10'd74  : rgb_data = 0;
10'd75  : rgb_data = 0;
10'd76  : rgb_data = 236;
10'd77  : rgb_data = 236;
10'd78  : rgb_data = 236;
10'd79  : rgb_data = 236;
10'd80  : rgb_data = 236;
10'd81  : rgb_data = 236;
10'd82  : rgb_data = 236;
10'd83  : rgb_data = 236;
10'd84  : rgb_data = 0;
10'd85  : rgb_data = 0;
10'd86  : rgb_data = 0;
10'd87  : rgb_data = 0;
10'd88  : rgb_data = 0;
10'd89  : rgb_data = 0;
10'd90  : rgb_data = 0;
10'd91  : rgb_data = 0;
10'd92  : rgb_data = 0;
10'd93  : rgb_data = 0;
10'd94  : rgb_data = 0;
10'd95  : rgb_data = 0;
10'd96  : rgb_data = 0;
10'd97  : rgb_data = 0;
10'd98  : rgb_data = 0;
10'd99  : rgb_data = 0;
10'd100 : rgb_data = 0;
10'd101 : rgb_data = 0;
10'd102 : rgb_data = 0;
10'd103 : rgb_data = 0;
10'd104 : rgb_data = 0;
10'd105 : rgb_data = 0;
10'd106 : rgb_data = 0;
10'd107 : rgb_data = 0;
10'd108 : rgb_data = 236;
10'd109 : rgb_data = 236;
10'd110 : rgb_data = 236;
10'd111 : rgb_data = 236;
10'd112 : rgb_data = 236;
10'd113 : rgb_data = 236;
10'd114 : rgb_data = 236;
10'd115 : rgb_data = 236;
10'd116 : rgb_data = 0;
10'd117 : rgb_data = 0;
10'd118 : rgb_data = 0;
10'd119 : rgb_data = 0;
10'd120 : rgb_data = 0;
10'd121 : rgb_data = 0;
10'd122 : rgb_data = 0;
10'd123 : rgb_data = 0;
10'd124 : rgb_data = 0;
10'd125 : rgb_data = 0;
10'd126 : rgb_data = 0;
10'd127 : rgb_data = 0;
10'd128 : rgb_data = 0;
10'd129 : rgb_data = 0;
10'd130 : rgb_data = 0;
10'd131 : rgb_data = 0;
10'd132 : rgb_data = 0;
10'd133 : rgb_data = 0;
10'd134 : rgb_data = 0;
10'd135 : rgb_data = 0;
10'd136 : rgb_data = 236;
10'd137 : rgb_data = 236;
10'd138 : rgb_data = 236;
10'd139 : rgb_data = 236;
10'd140 : rgb_data = 236;
10'd141 : rgb_data = 236;
10'd142 : rgb_data = 236;
10'd143 : rgb_data = 236;
10'd144 : rgb_data = 236;
10'd145 : rgb_data = 236;
10'd146 : rgb_data = 236;
10'd147 : rgb_data = 236;
10'd148 : rgb_data = 236;
10'd149 : rgb_data = 236;
10'd150 : rgb_data = 236;
10'd151 : rgb_data = 236;
10'd152 : rgb_data = 0;
10'd153 : rgb_data = 0;
10'd154 : rgb_data = 0;
10'd155 : rgb_data = 0;
10'd156 : rgb_data = 0;
10'd157 : rgb_data = 0;
10'd158 : rgb_data = 0;
10'd159 : rgb_data = 0;
10'd160 : rgb_data = 0;
10'd161 : rgb_data = 0;
10'd162 : rgb_data = 0;
10'd163 : rgb_data = 0;
10'd164 : rgb_data = 0;
10'd165 : rgb_data = 0;
10'd166 : rgb_data = 0;
10'd167 : rgb_data = 0;
10'd168 : rgb_data = 236;
10'd169 : rgb_data = 236;
10'd170 : rgb_data = 236;
10'd171 : rgb_data = 236;
10'd172 : rgb_data = 236;
10'd173 : rgb_data = 236;
10'd174 : rgb_data = 236;
10'd175 : rgb_data = 236;
10'd176 : rgb_data = 236;
10'd177 : rgb_data = 236;
10'd178 : rgb_data = 236;
10'd179 : rgb_data = 236;
10'd180 : rgb_data = 236;
10'd181 : rgb_data = 236;
10'd182 : rgb_data = 236;
10'd183 : rgb_data = 236;
10'd184 : rgb_data = 0;
10'd185 : rgb_data = 0;
10'd186 : rgb_data = 0;
10'd187 : rgb_data = 0;
10'd188 : rgb_data = 0;
10'd189 : rgb_data = 0;
10'd190 : rgb_data = 0;
10'd191 : rgb_data = 0;
10'd192 : rgb_data = 0;
10'd193 : rgb_data = 0;
10'd194 : rgb_data = 0;
10'd195 : rgb_data = 0;
10'd196 : rgb_data = 0;
10'd197 : rgb_data = 0;
10'd198 : rgb_data = 0;
10'd199 : rgb_data = 0;
10'd200 : rgb_data = 236;
10'd201 : rgb_data = 236;
10'd202 : rgb_data = 236;
10'd203 : rgb_data = 236;
10'd204 : rgb_data = 236;
10'd205 : rgb_data = 236;
10'd206 : rgb_data = 236;
10'd207 : rgb_data = 236;
10'd208 : rgb_data = 236;
10'd209 : rgb_data = 236;
10'd210 : rgb_data = 236;
10'd211 : rgb_data = 236;
10'd212 : rgb_data = 236;
10'd213 : rgb_data = 236;
10'd214 : rgb_data = 236;
10'd215 : rgb_data = 236;
10'd216 : rgb_data = 0;
10'd217 : rgb_data = 0;
10'd218 : rgb_data = 0;
10'd219 : rgb_data = 0;
10'd220 : rgb_data = 0;
10'd221 : rgb_data = 0;
10'd222 : rgb_data = 0;
10'd223 : rgb_data = 0;
10'd224 : rgb_data = 0;
10'd225 : rgb_data = 0;
10'd226 : rgb_data = 0;
10'd227 : rgb_data = 0;
10'd228 : rgb_data = 0;
10'd229 : rgb_data = 0;
10'd230 : rgb_data = 0;
10'd231 : rgb_data = 0;
10'd232 : rgb_data = 236;
10'd233 : rgb_data = 236;
10'd234 : rgb_data = 236;
10'd235 : rgb_data = 236;
10'd236 : rgb_data = 236;
10'd237 : rgb_data = 236;
10'd238 : rgb_data = 236;
10'd239 : rgb_data = 236;
10'd240 : rgb_data = 236;
10'd241 : rgb_data = 236;
10'd242 : rgb_data = 236;
10'd243 : rgb_data = 236;
10'd244 : rgb_data = 236;
10'd245 : rgb_data = 236;
10'd246 : rgb_data = 236;
10'd247 : rgb_data = 236;
10'd248 : rgb_data = 0;
10'd249 : rgb_data = 0;
10'd250 : rgb_data = 0;
10'd251 : rgb_data = 0;
10'd252 : rgb_data = 0;
10'd253 : rgb_data = 0;
10'd254 : rgb_data = 0;
10'd255 : rgb_data = 0;
10'd256 : rgb_data = 0;
10'd257 : rgb_data = 0;
10'd258 : rgb_data = 0;
10'd259 : rgb_data = 0;
10'd260 : rgb_data = 236;
10'd261 : rgb_data = 236;
10'd262 : rgb_data = 236;
10'd263 : rgb_data = 236;
10'd264 : rgb_data = 236;
10'd265 : rgb_data = 236;
10'd266 : rgb_data = 236;
10'd267 : rgb_data = 236;
10'd268 : rgb_data = 236;
10'd269 : rgb_data = 236;
10'd270 : rgb_data = 236;
10'd271 : rgb_data = 236;
10'd272 : rgb_data = 236;
10'd273 : rgb_data = 236;
10'd274 : rgb_data = 236;
10'd275 : rgb_data = 236;
10'd276 : rgb_data = 236;
10'd277 : rgb_data = 236;
10'd278 : rgb_data = 236;
10'd279 : rgb_data = 236;
10'd280 : rgb_data = 236;
10'd281 : rgb_data = 236;
10'd282 : rgb_data = 236;
10'd283 : rgb_data = 236;
10'd284 : rgb_data = 0;
10'd285 : rgb_data = 0;
10'd286 : rgb_data = 0;
10'd287 : rgb_data = 0;
10'd288 : rgb_data = 0;
10'd289 : rgb_data = 0;
10'd290 : rgb_data = 0;
10'd291 : rgb_data = 0;
10'd292 : rgb_data = 236;
10'd293 : rgb_data = 236;
10'd294 : rgb_data = 236;
10'd295 : rgb_data = 236;
10'd296 : rgb_data = 236;
10'd297 : rgb_data = 236;
10'd298 : rgb_data = 236;
10'd299 : rgb_data = 236;
10'd300 : rgb_data = 236;
10'd301 : rgb_data = 236;
10'd302 : rgb_data = 236;
10'd303 : rgb_data = 236;
10'd304 : rgb_data = 236;
10'd305 : rgb_data = 236;
10'd306 : rgb_data = 236;
10'd307 : rgb_data = 236;
10'd308 : rgb_data = 236;
10'd309 : rgb_data = 236;
10'd310 : rgb_data = 236;
10'd311 : rgb_data = 236;
10'd312 : rgb_data = 236;
10'd313 : rgb_data = 236;
10'd314 : rgb_data = 236;
10'd315 : rgb_data = 236;
10'd316 : rgb_data = 0;
10'd317 : rgb_data = 0;
10'd318 : rgb_data = 0;
10'd319 : rgb_data = 0;
10'd320 : rgb_data = 0;
10'd321 : rgb_data = 0;
10'd322 : rgb_data = 0;
10'd323 : rgb_data = 0;
10'd324 : rgb_data = 236;
10'd325 : rgb_data = 236;
10'd326 : rgb_data = 236;
10'd327 : rgb_data = 236;
10'd328 : rgb_data = 236;
10'd329 : rgb_data = 236;
10'd330 : rgb_data = 236;
10'd331 : rgb_data = 236;
10'd332 : rgb_data = 236;
10'd333 : rgb_data = 236;
10'd334 : rgb_data = 236;
10'd335 : rgb_data = 236;
10'd336 : rgb_data = 236;
10'd337 : rgb_data = 236;
10'd338 : rgb_data = 236;
10'd339 : rgb_data = 236;
10'd340 : rgb_data = 236;
10'd341 : rgb_data = 236;
10'd342 : rgb_data = 236;
10'd343 : rgb_data = 236;
10'd344 : rgb_data = 236;
10'd345 : rgb_data = 236;
10'd346 : rgb_data = 236;
10'd347 : rgb_data = 236;
10'd348 : rgb_data = 0;
10'd349 : rgb_data = 0;
10'd350 : rgb_data = 0;
10'd351 : rgb_data = 0;
10'd352 : rgb_data = 0;
10'd353 : rgb_data = 0;
10'd354 : rgb_data = 0;
10'd355 : rgb_data = 0;
10'd356 : rgb_data = 236;
10'd357 : rgb_data = 236;
10'd358 : rgb_data = 236;
10'd359 : rgb_data = 236;
10'd360 : rgb_data = 0;
10'd361 : rgb_data = 0;
10'd362 : rgb_data = 0;
10'd363 : rgb_data = 0;
10'd364 : rgb_data = 236;
10'd365 : rgb_data = 236;
10'd366 : rgb_data = 236;
10'd367 : rgb_data = 236;
10'd368 : rgb_data = 236;
10'd369 : rgb_data = 236;
10'd370 : rgb_data = 236;
10'd371 : rgb_data = 236;
10'd372 : rgb_data = 0;
10'd373 : rgb_data = 0;
10'd374 : rgb_data = 0;
10'd375 : rgb_data = 0;
10'd376 : rgb_data = 236;
10'd377 : rgb_data = 236;
10'd378 : rgb_data = 236;
10'd379 : rgb_data = 236;
10'd380 : rgb_data = 0;
10'd381 : rgb_data = 0;
10'd382 : rgb_data = 0;
10'd383 : rgb_data = 0;
10'd384 : rgb_data = 236;
10'd385 : rgb_data = 236;
10'd386 : rgb_data = 236;
10'd387 : rgb_data = 236;
10'd388 : rgb_data = 236;
10'd389 : rgb_data = 236;
10'd390 : rgb_data = 236;
10'd391 : rgb_data = 236;
10'd392 : rgb_data = 0;
10'd393 : rgb_data = 0;
10'd394 : rgb_data = 0;
10'd395 : rgb_data = 0;
10'd396 : rgb_data = 236;
10'd397 : rgb_data = 236;
10'd398 : rgb_data = 236;
10'd399 : rgb_data = 236;
10'd400 : rgb_data = 236;
10'd401 : rgb_data = 236;
10'd402 : rgb_data = 236;
10'd403 : rgb_data = 236;
10'd404 : rgb_data = 0;
10'd405 : rgb_data = 0;
10'd406 : rgb_data = 0;
10'd407 : rgb_data = 0;
10'd408 : rgb_data = 236;
10'd409 : rgb_data = 236;
10'd410 : rgb_data = 236;
10'd411 : rgb_data = 236;
10'd412 : rgb_data = 236;
10'd413 : rgb_data = 236;
10'd414 : rgb_data = 236;
10'd415 : rgb_data = 236;
10'd416 : rgb_data = 236;
10'd417 : rgb_data = 236;
10'd418 : rgb_data = 236;
10'd419 : rgb_data = 236;
10'd420 : rgb_data = 236;
10'd421 : rgb_data = 236;
10'd422 : rgb_data = 236;
10'd423 : rgb_data = 236;
10'd424 : rgb_data = 0;
10'd425 : rgb_data = 0;
10'd426 : rgb_data = 0;
10'd427 : rgb_data = 0;
10'd428 : rgb_data = 236;
10'd429 : rgb_data = 236;
10'd430 : rgb_data = 236;
10'd431 : rgb_data = 236;
10'd432 : rgb_data = 236;
10'd433 : rgb_data = 236;
10'd434 : rgb_data = 236;
10'd435 : rgb_data = 236;
10'd436 : rgb_data = 0;
10'd437 : rgb_data = 0;
10'd438 : rgb_data = 0;
10'd439 : rgb_data = 0;
10'd440 : rgb_data = 236;
10'd441 : rgb_data = 236;
10'd442 : rgb_data = 236;
10'd443 : rgb_data = 236;
10'd444 : rgb_data = 236;
10'd445 : rgb_data = 236;
10'd446 : rgb_data = 236;
10'd447 : rgb_data = 236;
10'd448 : rgb_data = 236;
10'd449 : rgb_data = 236;
10'd450 : rgb_data = 236;
10'd451 : rgb_data = 236;
10'd452 : rgb_data = 236;
10'd453 : rgb_data = 236;
10'd454 : rgb_data = 236;
10'd455 : rgb_data = 236;
10'd456 : rgb_data = 0;
10'd457 : rgb_data = 0;
10'd458 : rgb_data = 0;
10'd459 : rgb_data = 0;
10'd460 : rgb_data = 236;
10'd461 : rgb_data = 236;
10'd462 : rgb_data = 236;
10'd463 : rgb_data = 236;
10'd464 : rgb_data = 236;
10'd465 : rgb_data = 236;
10'd466 : rgb_data = 236;
10'd467 : rgb_data = 236;
10'd468 : rgb_data = 0;
10'd469 : rgb_data = 0;
10'd470 : rgb_data = 0;
10'd471 : rgb_data = 0;
10'd472 : rgb_data = 236;
10'd473 : rgb_data = 236;
10'd474 : rgb_data = 236;
10'd475 : rgb_data = 236;
10'd476 : rgb_data = 236;
10'd477 : rgb_data = 236;
10'd478 : rgb_data = 236;
10'd479 : rgb_data = 236;
10'd480 : rgb_data = 236;
10'd481 : rgb_data = 236;
10'd482 : rgb_data = 236;
10'd483 : rgb_data = 236;
10'd484 : rgb_data = 236;
10'd485 : rgb_data = 236;
10'd486 : rgb_data = 236;
10'd487 : rgb_data = 236;
10'd488 : rgb_data = 236;
10'd489 : rgb_data = 236;
10'd490 : rgb_data = 236;
10'd491 : rgb_data = 236;
10'd492 : rgb_data = 236;
10'd493 : rgb_data = 236;
10'd494 : rgb_data = 236;
10'd495 : rgb_data = 236;
10'd496 : rgb_data = 236;
10'd497 : rgb_data = 236;
10'd498 : rgb_data = 236;
10'd499 : rgb_data = 236;
10'd500 : rgb_data = 236;
10'd501 : rgb_data = 236;
10'd502 : rgb_data = 236;
10'd503 : rgb_data = 236;
10'd504 : rgb_data = 236;
10'd505 : rgb_data = 236;
10'd506 : rgb_data = 236;
10'd507 : rgb_data = 236;
10'd508 : rgb_data = 236;
10'd509 : rgb_data = 236;
10'd510 : rgb_data = 236;
10'd511 : rgb_data = 236;
10'd512 : rgb_data = 236;
10'd513 : rgb_data = 236;
10'd514 : rgb_data = 236;
10'd515 : rgb_data = 236;
10'd516 : rgb_data = 236;
10'd517 : rgb_data = 236;
10'd518 : rgb_data = 236;
10'd519 : rgb_data = 236;
10'd520 : rgb_data = 236;
10'd521 : rgb_data = 236;
10'd522 : rgb_data = 236;
10'd523 : rgb_data = 236;
10'd524 : rgb_data = 236;
10'd525 : rgb_data = 236;
10'd526 : rgb_data = 236;
10'd527 : rgb_data = 236;
10'd528 : rgb_data = 236;
10'd529 : rgb_data = 236;
10'd530 : rgb_data = 236;
10'd531 : rgb_data = 236;
10'd532 : rgb_data = 236;
10'd533 : rgb_data = 236;
10'd534 : rgb_data = 236;
10'd535 : rgb_data = 236;
10'd536 : rgb_data = 236;
10'd537 : rgb_data = 236;
10'd538 : rgb_data = 236;
10'd539 : rgb_data = 236;
10'd540 : rgb_data = 236;
10'd541 : rgb_data = 236;
10'd542 : rgb_data = 236;
10'd543 : rgb_data = 236;
10'd544 : rgb_data = 236;
10'd545 : rgb_data = 236;
10'd546 : rgb_data = 236;
10'd547 : rgb_data = 236;
10'd548 : rgb_data = 236;
10'd549 : rgb_data = 236;
10'd550 : rgb_data = 236;
10'd551 : rgb_data = 236;
10'd552 : rgb_data = 236;
10'd553 : rgb_data = 236;
10'd554 : rgb_data = 236;
10'd555 : rgb_data = 236;
10'd556 : rgb_data = 236;
10'd557 : rgb_data = 236;
10'd558 : rgb_data = 236;
10'd559 : rgb_data = 236;
10'd560 : rgb_data = 236;
10'd561 : rgb_data = 236;
10'd562 : rgb_data = 236;
10'd563 : rgb_data = 236;
10'd564 : rgb_data = 236;
10'd565 : rgb_data = 236;
10'd566 : rgb_data = 236;
10'd567 : rgb_data = 236;
10'd568 : rgb_data = 236;
10'd569 : rgb_data = 236;
10'd570 : rgb_data = 236;
10'd571 : rgb_data = 236;
10'd572 : rgb_data = 236;
10'd573 : rgb_data = 236;
10'd574 : rgb_data = 236;
10'd575 : rgb_data = 236;
10'd576 : rgb_data = 236;
10'd577 : rgb_data = 236;
10'd578 : rgb_data = 236;
10'd579 : rgb_data = 236;
10'd580 : rgb_data = 236;
10'd581 : rgb_data = 236;
10'd582 : rgb_data = 236;
10'd583 : rgb_data = 236;
10'd584 : rgb_data = 236;
10'd585 : rgb_data = 236;
10'd586 : rgb_data = 236;
10'd587 : rgb_data = 236;
10'd588 : rgb_data = 236;
10'd589 : rgb_data = 236;
10'd590 : rgb_data = 236;
10'd591 : rgb_data = 236;
10'd592 : rgb_data = 236;
10'd593 : rgb_data = 236;
10'd594 : rgb_data = 236;
10'd595 : rgb_data = 236;
10'd596 : rgb_data = 236;
10'd597 : rgb_data = 236;
10'd598 : rgb_data = 236;
10'd599 : rgb_data = 236;
10'd600 : rgb_data = 236;
10'd601 : rgb_data = 236;
10'd602 : rgb_data = 236;
10'd603 : rgb_data = 236;
10'd604 : rgb_data = 236;
10'd605 : rgb_data = 236;
10'd606 : rgb_data = 236;
10'd607 : rgb_data = 236;
10'd608 : rgb_data = 236;
10'd609 : rgb_data = 236;
10'd610 : rgb_data = 236;
10'd611 : rgb_data = 236;
10'd612 : rgb_data = 236;
10'd613 : rgb_data = 236;
10'd614 : rgb_data = 236;
10'd615 : rgb_data = 236;
10'd616 : rgb_data = 236;
10'd617 : rgb_data = 236;
10'd618 : rgb_data = 236;
10'd619 : rgb_data = 236;
10'd620 : rgb_data = 236;
10'd621 : rgb_data = 236;
10'd622 : rgb_data = 236;
10'd623 : rgb_data = 236;
10'd624 : rgb_data = 236;
10'd625 : rgb_data = 236;
10'd626 : rgb_data = 236;
10'd627 : rgb_data = 236;
10'd628 : rgb_data = 236;
10'd629 : rgb_data = 236;
10'd630 : rgb_data = 236;
10'd631 : rgb_data = 236;
10'd632 : rgb_data = 236;
10'd633 : rgb_data = 236;
10'd634 : rgb_data = 236;
10'd635 : rgb_data = 236;
10'd636 : rgb_data = 236;
10'd637 : rgb_data = 236;
10'd638 : rgb_data = 236;
10'd639 : rgb_data = 236;
10'd640 : rgb_data = 0;
10'd641 : rgb_data = 0;
10'd642 : rgb_data = 0;
10'd643 : rgb_data = 0;
10'd644 : rgb_data = 0;
10'd645 : rgb_data = 0;
10'd646 : rgb_data = 0;
10'd647 : rgb_data = 0;
10'd648 : rgb_data = 236;
10'd649 : rgb_data = 236;
10'd650 : rgb_data = 236;
10'd651 : rgb_data = 236;
10'd652 : rgb_data = 0;
10'd653 : rgb_data = 0;
10'd654 : rgb_data = 0;
10'd655 : rgb_data = 0;
10'd656 : rgb_data = 0;
10'd657 : rgb_data = 0;
10'd658 : rgb_data = 0;
10'd659 : rgb_data = 0;
10'd660 : rgb_data = 236;
10'd661 : rgb_data = 236;
10'd662 : rgb_data = 236;
10'd663 : rgb_data = 236;
10'd664 : rgb_data = 0;
10'd665 : rgb_data = 0;
10'd666 : rgb_data = 0;
10'd667 : rgb_data = 0;
10'd668 : rgb_data = 0;
10'd669 : rgb_data = 0;
10'd670 : rgb_data = 0;
10'd671 : rgb_data = 0;
10'd672 : rgb_data = 0;
10'd673 : rgb_data = 0;
10'd674 : rgb_data = 0;
10'd675 : rgb_data = 0;
10'd676 : rgb_data = 0;
10'd677 : rgb_data = 0;
10'd678 : rgb_data = 0;
10'd679 : rgb_data = 0;
10'd680 : rgb_data = 236;
10'd681 : rgb_data = 236;
10'd682 : rgb_data = 236;
10'd683 : rgb_data = 236;
10'd684 : rgb_data = 0;
10'd685 : rgb_data = 0;
10'd686 : rgb_data = 0;
10'd687 : rgb_data = 0;
10'd688 : rgb_data = 0;
10'd689 : rgb_data = 0;
10'd690 : rgb_data = 0;
10'd691 : rgb_data = 0;
10'd692 : rgb_data = 236;
10'd693 : rgb_data = 236;
10'd694 : rgb_data = 236;
10'd695 : rgb_data = 236;
10'd696 : rgb_data = 0;
10'd697 : rgb_data = 0;
10'd698 : rgb_data = 0;
10'd699 : rgb_data = 0;
10'd700 : rgb_data = 0;
10'd701 : rgb_data = 0;
10'd702 : rgb_data = 0;
10'd703 : rgb_data = 0;
10'd704 : rgb_data = 0;
10'd705 : rgb_data = 0;
10'd706 : rgb_data = 0;
10'd707 : rgb_data = 0;
10'd708 : rgb_data = 0;
10'd709 : rgb_data = 0;
10'd710 : rgb_data = 0;
10'd711 : rgb_data = 0;
10'd712 : rgb_data = 236;
10'd713 : rgb_data = 236;
10'd714 : rgb_data = 236;
10'd715 : rgb_data = 236;
10'd716 : rgb_data = 0;
10'd717 : rgb_data = 0;
10'd718 : rgb_data = 0;
10'd719 : rgb_data = 0;
10'd720 : rgb_data = 0;
10'd721 : rgb_data = 0;
10'd722 : rgb_data = 0;
10'd723 : rgb_data = 0;
10'd724 : rgb_data = 236;
10'd725 : rgb_data = 236;
10'd726 : rgb_data = 236;
10'd727 : rgb_data = 236;
10'd728 : rgb_data = 0;
10'd729 : rgb_data = 0;
10'd730 : rgb_data = 0;
10'd731 : rgb_data = 0;
10'd732 : rgb_data = 0;
10'd733 : rgb_data = 0;
10'd734 : rgb_data = 0;
10'd735 : rgb_data = 0;
10'd736 : rgb_data = 0;
10'd737 : rgb_data = 0;
10'd738 : rgb_data = 0;
10'd739 : rgb_data = 0;
10'd740 : rgb_data = 0;
10'd741 : rgb_data = 0;
10'd742 : rgb_data = 0;
10'd743 : rgb_data = 0;
10'd744 : rgb_data = 236;
10'd745 : rgb_data = 236;
10'd746 : rgb_data = 236;
10'd747 : rgb_data = 236;
10'd748 : rgb_data = 0;
10'd749 : rgb_data = 0;
10'd750 : rgb_data = 0;
10'd751 : rgb_data = 0;
10'd752 : rgb_data = 0;
10'd753 : rgb_data = 0;
10'd754 : rgb_data = 0;
10'd755 : rgb_data = 0;
10'd756 : rgb_data = 236;
10'd757 : rgb_data = 236;
10'd758 : rgb_data = 236;
10'd759 : rgb_data = 236;
10'd760 : rgb_data = 0;
10'd761 : rgb_data = 0;
10'd762 : rgb_data = 0;
10'd763 : rgb_data = 0;
10'd764 : rgb_data = 0;
10'd765 : rgb_data = 0;
10'd766 : rgb_data = 0;
10'd767 : rgb_data = 0;
10'd768 : rgb_data = 0;
10'd769 : rgb_data = 0;
10'd770 : rgb_data = 0;
10'd771 : rgb_data = 0;
10'd772 : rgb_data = 236;
10'd773 : rgb_data = 236;
10'd774 : rgb_data = 236;
10'd775 : rgb_data = 236;
10'd776 : rgb_data = 0;
10'd777 : rgb_data = 0;
10'd778 : rgb_data = 0;
10'd779 : rgb_data = 0;
10'd780 : rgb_data = 236;
10'd781 : rgb_data = 236;
10'd782 : rgb_data = 236;
10'd783 : rgb_data = 236;
10'd784 : rgb_data = 236;
10'd785 : rgb_data = 236;
10'd786 : rgb_data = 236;
10'd787 : rgb_data = 236;
10'd788 : rgb_data = 0;
10'd789 : rgb_data = 0;
10'd790 : rgb_data = 0;
10'd791 : rgb_data = 0;
10'd792 : rgb_data = 236;
10'd793 : rgb_data = 236;
10'd794 : rgb_data = 236;
10'd795 : rgb_data = 236;
10'd796 : rgb_data = 0;
10'd797 : rgb_data = 0;
10'd798 : rgb_data = 0;
10'd799 : rgb_data = 0;
10'd800 : rgb_data = 0;
10'd801 : rgb_data = 0;
10'd802 : rgb_data = 0;
10'd803 : rgb_data = 0;
10'd804 : rgb_data = 236;
10'd805 : rgb_data = 236;
10'd806 : rgb_data = 236;
10'd807 : rgb_data = 236;
10'd808 : rgb_data = 0;
10'd809 : rgb_data = 0;
10'd810 : rgb_data = 0;
10'd811 : rgb_data = 0;
10'd812 : rgb_data = 236;
10'd813 : rgb_data = 236;
10'd814 : rgb_data = 236;
10'd815 : rgb_data = 236;
10'd816 : rgb_data = 236;
10'd817 : rgb_data = 236;
10'd818 : rgb_data = 236;
10'd819 : rgb_data = 236;
10'd820 : rgb_data = 0;
10'd821 : rgb_data = 0;
10'd822 : rgb_data = 0;
10'd823 : rgb_data = 0;
10'd824 : rgb_data = 236;
10'd825 : rgb_data = 236;
10'd826 : rgb_data = 236;
10'd827 : rgb_data = 236;
10'd828 : rgb_data = 0;
10'd829 : rgb_data = 0;
10'd830 : rgb_data = 0;
10'd831 : rgb_data = 0;
10'd832 : rgb_data = 0;
10'd833 : rgb_data = 0;
10'd834 : rgb_data = 0;
10'd835 : rgb_data = 0;
10'd836 : rgb_data = 236;
10'd837 : rgb_data = 236;
10'd838 : rgb_data = 236;
10'd839 : rgb_data = 236;
10'd840 : rgb_data = 0;
10'd841 : rgb_data = 0;
10'd842 : rgb_data = 0;
10'd843 : rgb_data = 0;
10'd844 : rgb_data = 236;
10'd845 : rgb_data = 236;
10'd846 : rgb_data = 236;
10'd847 : rgb_data = 236;
10'd848 : rgb_data = 236;
10'd849 : rgb_data = 236;
10'd850 : rgb_data = 236;
10'd851 : rgb_data = 236;
10'd852 : rgb_data = 0;
10'd853 : rgb_data = 0;
10'd854 : rgb_data = 0;
10'd855 : rgb_data = 0;
10'd856 : rgb_data = 236;
10'd857 : rgb_data = 236;
10'd858 : rgb_data = 236;
10'd859 : rgb_data = 236;
10'd860 : rgb_data = 0;
10'd861 : rgb_data = 0;
10'd862 : rgb_data = 0;
10'd863 : rgb_data = 0;
10'd864 : rgb_data = 0;
10'd865 : rgb_data = 0;
10'd866 : rgb_data = 0;
10'd867 : rgb_data = 0;
10'd868 : rgb_data = 236;
10'd869 : rgb_data = 236;
10'd870 : rgb_data = 236;
10'd871 : rgb_data = 236;
10'd872 : rgb_data = 0;
10'd873 : rgb_data = 0;
10'd874 : rgb_data = 0;
10'd875 : rgb_data = 0;
10'd876 : rgb_data = 236;
10'd877 : rgb_data = 236;
10'd878 : rgb_data = 236;
10'd879 : rgb_data = 236;
10'd880 : rgb_data = 236;
10'd881 : rgb_data = 236;
10'd882 : rgb_data = 236;
10'd883 : rgb_data = 236;
10'd884 : rgb_data = 0;
10'd885 : rgb_data = 0;
10'd886 : rgb_data = 0;
10'd887 : rgb_data = 0;
10'd888 : rgb_data = 236;
10'd889 : rgb_data = 236;
10'd890 : rgb_data = 236;
10'd891 : rgb_data = 236;
10'd892 : rgb_data = 0;
10'd893 : rgb_data = 0;
10'd894 : rgb_data = 0;
10'd895 : rgb_data = 0;
10'd896 : rgb_data = 236;
10'd897 : rgb_data = 236;
10'd898 : rgb_data = 236;
10'd899 : rgb_data = 236;
10'd900 : rgb_data = 0;
10'd901 : rgb_data = 0;
10'd902 : rgb_data = 0;
10'd903 : rgb_data = 0;
10'd904 : rgb_data = 236;
10'd905 : rgb_data = 236;
10'd906 : rgb_data = 236;
10'd907 : rgb_data = 236;
10'd908 : rgb_data = 0;
10'd909 : rgb_data = 0;
10'd910 : rgb_data = 0;
10'd911 : rgb_data = 0;
10'd912 : rgb_data = 0;
10'd913 : rgb_data = 0;
10'd914 : rgb_data = 0;
10'd915 : rgb_data = 0;
10'd916 : rgb_data = 236;
10'd917 : rgb_data = 236;
10'd918 : rgb_data = 236;
10'd919 : rgb_data = 236;
10'd920 : rgb_data = 0;
10'd921 : rgb_data = 0;
10'd922 : rgb_data = 0;
10'd923 : rgb_data = 0;
10'd924 : rgb_data = 236;
10'd925 : rgb_data = 236;
10'd926 : rgb_data = 236;
10'd927 : rgb_data = 236;
10'd928 : rgb_data = 236;
10'd929 : rgb_data = 236;
10'd930 : rgb_data = 236;
10'd931 : rgb_data = 236;
10'd932 : rgb_data = 0;
10'd933 : rgb_data = 0;
10'd934 : rgb_data = 0;
10'd935 : rgb_data = 0;
10'd936 : rgb_data = 236;
10'd937 : rgb_data = 236;
10'd938 : rgb_data = 236;
10'd939 : rgb_data = 236;
10'd940 : rgb_data = 0;
10'd941 : rgb_data = 0;
10'd942 : rgb_data = 0;
10'd943 : rgb_data = 0;
10'd944 : rgb_data = 0;
10'd945 : rgb_data = 0;
10'd946 : rgb_data = 0;
10'd947 : rgb_data = 0;
10'd948 : rgb_data = 236;
10'd949 : rgb_data = 236;
10'd950 : rgb_data = 236;
10'd951 : rgb_data = 236;
10'd952 : rgb_data = 0;
10'd953 : rgb_data = 0;
10'd954 : rgb_data = 0;
10'd955 : rgb_data = 0;
10'd956 : rgb_data = 236;
10'd957 : rgb_data = 236;
10'd958 : rgb_data = 236;
10'd959 : rgb_data = 236;
10'd960 : rgb_data = 236;
10'd961 : rgb_data = 236;
10'd962 : rgb_data = 236;
10'd963 : rgb_data = 236;
10'd964 : rgb_data = 0;
10'd965 : rgb_data = 0;
10'd966 : rgb_data = 0;
10'd967 : rgb_data = 0;
10'd968 : rgb_data = 236;
10'd969 : rgb_data = 236;
10'd970 : rgb_data = 236;
10'd971 : rgb_data = 236;
10'd972 : rgb_data = 0;
10'd973 : rgb_data = 0;
10'd974 : rgb_data = 0;
10'd975 : rgb_data = 0;
10'd976 : rgb_data = 0;
10'd977 : rgb_data = 0;
10'd978 : rgb_data = 0;
10'd979 : rgb_data = 0;
10'd980 : rgb_data = 236;
10'd981 : rgb_data = 236;
10'd982 : rgb_data = 236;
10'd983 : rgb_data = 236;
10'd984 : rgb_data = 0;
10'd985 : rgb_data = 0;
10'd986 : rgb_data = 0;
10'd987 : rgb_data = 0;
10'd988 : rgb_data = 236;
10'd989 : rgb_data = 236;
10'd990 : rgb_data = 236;
10'd991 : rgb_data = 236;
10'd992 : rgb_data = 236;
10'd993 : rgb_data = 236;
10'd994 : rgb_data = 236;
10'd995 : rgb_data = 236;
10'd996 : rgb_data = 0;
10'd997 : rgb_data = 0;
10'd998 : rgb_data = 0;
10'd999 : rgb_data = 0;
10'd1000: rgb_data = 236;
10'd1001: rgb_data = 236;
10'd1002: rgb_data = 236;
10'd1003: rgb_data = 236;
10'd1004: rgb_data = 0;
10'd1005: rgb_data = 0;
10'd1006: rgb_data = 0;
10'd1007: rgb_data = 0;
10'd1008: rgb_data = 0;
10'd1009: rgb_data = 0;
10'd1010: rgb_data = 0;
10'd1011: rgb_data = 0;
10'd1012: rgb_data = 236;
10'd1013: rgb_data = 236;
10'd1014: rgb_data = 236;
10'd1015: rgb_data = 236;
10'd1016: rgb_data = 0;
10'd1017: rgb_data = 0;
10'd1018: rgb_data = 0;
10'd1019: rgb_data = 0;
10'd1020: rgb_data = 236;
10'd1021: rgb_data = 236;
10'd1022: rgb_data = 236;
10'd1023: rgb_data = 236;

default : rgb_data = 8'd0;
endcase

endmodule
