`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:15:18 11/13/2018 
// Design Name: 
// Module Name:    ship_rom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ship_rom(
input [11:0] address,
output reg [7:0] rgb_data
    );
(* rom_style = "block" *)


always @*
case(address)
12'd0   : rgb_data = 0;
12'd1   : rgb_data = 0;
12'd2   : rgb_data = 0;
12'd3   : rgb_data = 0;
12'd4   : rgb_data = 0;
12'd5   : rgb_data = 0;
12'd6   : rgb_data = 0;
12'd7   : rgb_data = 0;
12'd8   : rgb_data = 0;
12'd9   : rgb_data = 0;
12'd10  : rgb_data = 0;
12'd11  : rgb_data = 0;
12'd12  : rgb_data = 0;
12'd13  : rgb_data = 0;
12'd14  : rgb_data = 0;
12'd15  : rgb_data = 0;
12'd16  : rgb_data = 0;
12'd17  : rgb_data = 0;
12'd18  : rgb_data = 0;
12'd19  : rgb_data = 0;
12'd20  : rgb_data = 0;
12'd21  : rgb_data = 0;
12'd22  : rgb_data = 0;
12'd23  : rgb_data = 0;
12'd24  : rgb_data = 0;
12'd25  : rgb_data = 0;
12'd26  : rgb_data = 0;
12'd27  : rgb_data = 0;
12'd28  : rgb_data = 20;
12'd29  : rgb_data = 20;
12'd30  : rgb_data = 20;
12'd31  : rgb_data = 20;
12'd32  : rgb_data = 20;
12'd33  : rgb_data = 20;
12'd34  : rgb_data = 20;
12'd35  : rgb_data = 20;
12'd36  : rgb_data = 0;
12'd37  : rgb_data = 0;
12'd38  : rgb_data = 0;
12'd39  : rgb_data = 0;
12'd40  : rgb_data = 0;
12'd41  : rgb_data = 0;
12'd42  : rgb_data = 0;
12'd43  : rgb_data = 0;
12'd44  : rgb_data = 0;
12'd45  : rgb_data = 0;
12'd46  : rgb_data = 0;
12'd47  : rgb_data = 0;
12'd48  : rgb_data = 0;
12'd49  : rgb_data = 0;
12'd50  : rgb_data = 0;
12'd51  : rgb_data = 0;
12'd52  : rgb_data = 0;
12'd53  : rgb_data = 0;
12'd54  : rgb_data = 0;
12'd55  : rgb_data = 0;
12'd56  : rgb_data = 0;
12'd57  : rgb_data = 0;
12'd58  : rgb_data = 0;
12'd59  : rgb_data = 0;
12'd60  : rgb_data = 0;
12'd61  : rgb_data = 0;
12'd62  : rgb_data = 0;
12'd63  : rgb_data = 0;
12'd64  : rgb_data = 0;
12'd65  : rgb_data = 0;
12'd66  : rgb_data = 0;
12'd67  : rgb_data = 0;
12'd68  : rgb_data = 0;
12'd69  : rgb_data = 0;
12'd70  : rgb_data = 0;
12'd71  : rgb_data = 0;
12'd72  : rgb_data = 0;
12'd73  : rgb_data = 0;
12'd74  : rgb_data = 0;
12'd75  : rgb_data = 0;
12'd76  : rgb_data = 0;
12'd77  : rgb_data = 0;
12'd78  : rgb_data = 0;
12'd79  : rgb_data = 0;
12'd80  : rgb_data = 0;
12'd81  : rgb_data = 0;
12'd82  : rgb_data = 0;
12'd83  : rgb_data = 0;
12'd84  : rgb_data = 0;
12'd85  : rgb_data = 0;
12'd86  : rgb_data = 0;
12'd87  : rgb_data = 0;
12'd88  : rgb_data = 0;
12'd89  : rgb_data = 0;
12'd90  : rgb_data = 0;
12'd91  : rgb_data = 0;
12'd92  : rgb_data = 20;
12'd93  : rgb_data = 20;
12'd94  : rgb_data = 20;
12'd95  : rgb_data = 20;
12'd96  : rgb_data = 20;
12'd97  : rgb_data = 20;
12'd98  : rgb_data = 20;
12'd99  : rgb_data = 20;
12'd100 : rgb_data = 0;
12'd101 : rgb_data = 0;
12'd102 : rgb_data = 0;
12'd103 : rgb_data = 0;
12'd104 : rgb_data = 0;
12'd105 : rgb_data = 0;
12'd106 : rgb_data = 0;
12'd107 : rgb_data = 0;
12'd108 : rgb_data = 0;
12'd109 : rgb_data = 0;
12'd110 : rgb_data = 0;
12'd111 : rgb_data = 0;
12'd112 : rgb_data = 0;
12'd113 : rgb_data = 0;
12'd114 : rgb_data = 0;
12'd115 : rgb_data = 0;
12'd116 : rgb_data = 0;
12'd117 : rgb_data = 0;
12'd118 : rgb_data = 0;
12'd119 : rgb_data = 0;
12'd120 : rgb_data = 0;
12'd121 : rgb_data = 0;
12'd122 : rgb_data = 0;
12'd123 : rgb_data = 0;
12'd124 : rgb_data = 0;
12'd125 : rgb_data = 0;
12'd126 : rgb_data = 0;
12'd127 : rgb_data = 0;
12'd128 : rgb_data = 0;
12'd129 : rgb_data = 0;
12'd130 : rgb_data = 0;
12'd131 : rgb_data = 0;
12'd132 : rgb_data = 0;
12'd133 : rgb_data = 0;
12'd134 : rgb_data = 0;
12'd135 : rgb_data = 0;
12'd136 : rgb_data = 0;
12'd137 : rgb_data = 0;
12'd138 : rgb_data = 0;
12'd139 : rgb_data = 0;
12'd140 : rgb_data = 0;
12'd141 : rgb_data = 0;
12'd142 : rgb_data = 0;
12'd143 : rgb_data = 0;
12'd144 : rgb_data = 0;
12'd145 : rgb_data = 0;
12'd146 : rgb_data = 0;
12'd147 : rgb_data = 0;
12'd148 : rgb_data = 0;
12'd149 : rgb_data = 0;
12'd150 : rgb_data = 0;
12'd151 : rgb_data = 0;
12'd152 : rgb_data = 0;
12'd153 : rgb_data = 0;
12'd154 : rgb_data = 0;
12'd155 : rgb_data = 0;
12'd156 : rgb_data = 255;
12'd157 : rgb_data = 255;
12'd158 : rgb_data = 255;
12'd159 : rgb_data = 255;
12'd160 : rgb_data = 255;
12'd161 : rgb_data = 255;
12'd162 : rgb_data = 255;
12'd163 : rgb_data = 255;
12'd164 : rgb_data = 0;
12'd165 : rgb_data = 0;
12'd166 : rgb_data = 0;
12'd167 : rgb_data = 0;
12'd168 : rgb_data = 0;
12'd169 : rgb_data = 0;
12'd170 : rgb_data = 0;
12'd171 : rgb_data = 0;
12'd172 : rgb_data = 0;
12'd173 : rgb_data = 0;
12'd174 : rgb_data = 0;
12'd175 : rgb_data = 0;
12'd176 : rgb_data = 0;
12'd177 : rgb_data = 0;
12'd178 : rgb_data = 0;
12'd179 : rgb_data = 0;
12'd180 : rgb_data = 0;
12'd181 : rgb_data = 0;
12'd182 : rgb_data = 0;
12'd183 : rgb_data = 0;
12'd184 : rgb_data = 0;
12'd185 : rgb_data = 0;
12'd186 : rgb_data = 0;
12'd187 : rgb_data = 0;
12'd188 : rgb_data = 0;
12'd189 : rgb_data = 0;
12'd190 : rgb_data = 0;
12'd191 : rgb_data = 0;
12'd192 : rgb_data = 0;
12'd193 : rgb_data = 0;
12'd194 : rgb_data = 0;
12'd195 : rgb_data = 0;
12'd196 : rgb_data = 0;
12'd197 : rgb_data = 0;
12'd198 : rgb_data = 0;
12'd199 : rgb_data = 0;
12'd200 : rgb_data = 0;
12'd201 : rgb_data = 0;
12'd202 : rgb_data = 0;
12'd203 : rgb_data = 0;
12'd204 : rgb_data = 0;
12'd205 : rgb_data = 0;
12'd206 : rgb_data = 0;
12'd207 : rgb_data = 0;
12'd208 : rgb_data = 0;
12'd209 : rgb_data = 0;
12'd210 : rgb_data = 0;
12'd211 : rgb_data = 0;
12'd212 : rgb_data = 0;
12'd213 : rgb_data = 0;
12'd214 : rgb_data = 0;
12'd215 : rgb_data = 0;
12'd216 : rgb_data = 0;
12'd217 : rgb_data = 0;
12'd218 : rgb_data = 0;
12'd219 : rgb_data = 0;
12'd220 : rgb_data = 255;
12'd221 : rgb_data = 255;
12'd222 : rgb_data = 255;
12'd223 : rgb_data = 255;
12'd224 : rgb_data = 255;
12'd225 : rgb_data = 255;
12'd226 : rgb_data = 255;
12'd227 : rgb_data = 255;
12'd228 : rgb_data = 0;
12'd229 : rgb_data = 0;
12'd230 : rgb_data = 0;
12'd231 : rgb_data = 0;
12'd232 : rgb_data = 0;
12'd233 : rgb_data = 0;
12'd234 : rgb_data = 0;
12'd235 : rgb_data = 0;
12'd236 : rgb_data = 0;
12'd237 : rgb_data = 0;
12'd238 : rgb_data = 0;
12'd239 : rgb_data = 0;
12'd240 : rgb_data = 0;
12'd241 : rgb_data = 0;
12'd242 : rgb_data = 0;
12'd243 : rgb_data = 0;
12'd244 : rgb_data = 0;
12'd245 : rgb_data = 0;
12'd246 : rgb_data = 0;
12'd247 : rgb_data = 0;
12'd248 : rgb_data = 0;
12'd249 : rgb_data = 0;
12'd250 : rgb_data = 0;
12'd251 : rgb_data = 0;
12'd252 : rgb_data = 0;
12'd253 : rgb_data = 0;
12'd254 : rgb_data = 0;
12'd255 : rgb_data = 0;
12'd256 : rgb_data = 0;
12'd257 : rgb_data = 0;
12'd258 : rgb_data = 0;
12'd259 : rgb_data = 0;
12'd260 : rgb_data = 0;
12'd261 : rgb_data = 0;
12'd262 : rgb_data = 0;
12'd263 : rgb_data = 0;
12'd264 : rgb_data = 0;
12'd265 : rgb_data = 0;
12'd266 : rgb_data = 0;
12'd267 : rgb_data = 0;
12'd268 : rgb_data = 0;
12'd269 : rgb_data = 0;
12'd270 : rgb_data = 0;
12'd271 : rgb_data = 0;
12'd272 : rgb_data = 0;
12'd273 : rgb_data = 0;
12'd274 : rgb_data = 0;
12'd275 : rgb_data = 0;
12'd276 : rgb_data = 0;
12'd277 : rgb_data = 0;
12'd278 : rgb_data = 0;
12'd279 : rgb_data = 0;
12'd280 : rgb_data = 0;
12'd281 : rgb_data = 0;
12'd282 : rgb_data = 0;
12'd283 : rgb_data = 0;
12'd284 : rgb_data = 255;
12'd285 : rgb_data = 255;
12'd286 : rgb_data = 255;
12'd287 : rgb_data = 255;
12'd288 : rgb_data = 255;
12'd289 : rgb_data = 255;
12'd290 : rgb_data = 255;
12'd291 : rgb_data = 255;
12'd292 : rgb_data = 0;
12'd293 : rgb_data = 0;
12'd294 : rgb_data = 0;
12'd295 : rgb_data = 0;
12'd296 : rgb_data = 0;
12'd297 : rgb_data = 0;
12'd298 : rgb_data = 0;
12'd299 : rgb_data = 0;
12'd300 : rgb_data = 0;
12'd301 : rgb_data = 0;
12'd302 : rgb_data = 0;
12'd303 : rgb_data = 0;
12'd304 : rgb_data = 0;
12'd305 : rgb_data = 0;
12'd306 : rgb_data = 0;
12'd307 : rgb_data = 0;
12'd308 : rgb_data = 0;
12'd309 : rgb_data = 0;
12'd310 : rgb_data = 0;
12'd311 : rgb_data = 0;
12'd312 : rgb_data = 0;
12'd313 : rgb_data = 0;
12'd314 : rgb_data = 0;
12'd315 : rgb_data = 0;
12'd316 : rgb_data = 0;
12'd317 : rgb_data = 0;
12'd318 : rgb_data = 0;
12'd319 : rgb_data = 0;
12'd320 : rgb_data = 0;
12'd321 : rgb_data = 0;
12'd322 : rgb_data = 0;
12'd323 : rgb_data = 0;
12'd324 : rgb_data = 0;
12'd325 : rgb_data = 0;
12'd326 : rgb_data = 0;
12'd327 : rgb_data = 0;
12'd328 : rgb_data = 0;
12'd329 : rgb_data = 0;
12'd330 : rgb_data = 0;
12'd331 : rgb_data = 0;
12'd332 : rgb_data = 0;
12'd333 : rgb_data = 0;
12'd334 : rgb_data = 0;
12'd335 : rgb_data = 0;
12'd336 : rgb_data = 0;
12'd337 : rgb_data = 0;
12'd338 : rgb_data = 0;
12'd339 : rgb_data = 0;
12'd340 : rgb_data = 0;
12'd341 : rgb_data = 0;
12'd342 : rgb_data = 0;
12'd343 : rgb_data = 0;
12'd344 : rgb_data = 0;
12'd345 : rgb_data = 0;
12'd346 : rgb_data = 0;
12'd347 : rgb_data = 0;
12'd348 : rgb_data = 255;
12'd349 : rgb_data = 255;
12'd350 : rgb_data = 255;
12'd351 : rgb_data = 255;
12'd352 : rgb_data = 255;
12'd353 : rgb_data = 255;
12'd354 : rgb_data = 255;
12'd355 : rgb_data = 255;
12'd356 : rgb_data = 0;
12'd357 : rgb_data = 0;
12'd358 : rgb_data = 0;
12'd359 : rgb_data = 0;
12'd360 : rgb_data = 0;
12'd361 : rgb_data = 0;
12'd362 : rgb_data = 0;
12'd363 : rgb_data = 0;
12'd364 : rgb_data = 0;
12'd365 : rgb_data = 0;
12'd366 : rgb_data = 0;
12'd367 : rgb_data = 0;
12'd368 : rgb_data = 0;
12'd369 : rgb_data = 0;
12'd370 : rgb_data = 0;
12'd371 : rgb_data = 0;
12'd372 : rgb_data = 0;
12'd373 : rgb_data = 0;
12'd374 : rgb_data = 0;
12'd375 : rgb_data = 0;
12'd376 : rgb_data = 0;
12'd377 : rgb_data = 0;
12'd378 : rgb_data = 0;
12'd379 : rgb_data = 0;
12'd380 : rgb_data = 0;
12'd381 : rgb_data = 0;
12'd382 : rgb_data = 0;
12'd383 : rgb_data = 0;
12'd384 : rgb_data = 0;
12'd385 : rgb_data = 0;
12'd386 : rgb_data = 0;
12'd387 : rgb_data = 0;
12'd388 : rgb_data = 0;
12'd389 : rgb_data = 0;
12'd390 : rgb_data = 0;
12'd391 : rgb_data = 0;
12'd392 : rgb_data = 0;
12'd393 : rgb_data = 0;
12'd394 : rgb_data = 0;
12'd395 : rgb_data = 0;
12'd396 : rgb_data = 0;
12'd397 : rgb_data = 0;
12'd398 : rgb_data = 0;
12'd399 : rgb_data = 0;
12'd400 : rgb_data = 0;
12'd401 : rgb_data = 0;
12'd402 : rgb_data = 0;
12'd403 : rgb_data = 0;
12'd404 : rgb_data = 0;
12'd405 : rgb_data = 0;
12'd406 : rgb_data = 0;
12'd407 : rgb_data = 0;
12'd408 : rgb_data = 0;
12'd409 : rgb_data = 0;
12'd410 : rgb_data = 0;
12'd411 : rgb_data = 0;
12'd412 : rgb_data = 255;
12'd413 : rgb_data = 255;
12'd414 : rgb_data = 255;
12'd415 : rgb_data = 255;
12'd416 : rgb_data = 255;
12'd417 : rgb_data = 255;
12'd418 : rgb_data = 255;
12'd419 : rgb_data = 255;
12'd420 : rgb_data = 0;
12'd421 : rgb_data = 0;
12'd422 : rgb_data = 0;
12'd423 : rgb_data = 0;
12'd424 : rgb_data = 0;
12'd425 : rgb_data = 0;
12'd426 : rgb_data = 0;
12'd427 : rgb_data = 0;
12'd428 : rgb_data = 0;
12'd429 : rgb_data = 0;
12'd430 : rgb_data = 0;
12'd431 : rgb_data = 0;
12'd432 : rgb_data = 0;
12'd433 : rgb_data = 0;
12'd434 : rgb_data = 0;
12'd435 : rgb_data = 0;
12'd436 : rgb_data = 0;
12'd437 : rgb_data = 0;
12'd438 : rgb_data = 0;
12'd439 : rgb_data = 0;
12'd440 : rgb_data = 0;
12'd441 : rgb_data = 0;
12'd442 : rgb_data = 0;
12'd443 : rgb_data = 0;
12'd444 : rgb_data = 0;
12'd445 : rgb_data = 0;
12'd446 : rgb_data = 0;
12'd447 : rgb_data = 0;
12'd448 : rgb_data = 0;
12'd449 : rgb_data = 0;
12'd450 : rgb_data = 0;
12'd451 : rgb_data = 0;
12'd452 : rgb_data = 0;
12'd453 : rgb_data = 0;
12'd454 : rgb_data = 0;
12'd455 : rgb_data = 0;
12'd456 : rgb_data = 0;
12'd457 : rgb_data = 0;
12'd458 : rgb_data = 0;
12'd459 : rgb_data = 0;
12'd460 : rgb_data = 0;
12'd461 : rgb_data = 0;
12'd462 : rgb_data = 0;
12'd463 : rgb_data = 0;
12'd464 : rgb_data = 0;
12'd465 : rgb_data = 0;
12'd466 : rgb_data = 0;
12'd467 : rgb_data = 0;
12'd468 : rgb_data = 0;
12'd469 : rgb_data = 0;
12'd470 : rgb_data = 0;
12'd471 : rgb_data = 0;
12'd472 : rgb_data = 0;
12'd473 : rgb_data = 0;
12'd474 : rgb_data = 0;
12'd475 : rgb_data = 0;
12'd476 : rgb_data = 255;
12'd477 : rgb_data = 255;
12'd478 : rgb_data = 255;
12'd479 : rgb_data = 255;
12'd480 : rgb_data = 255;
12'd481 : rgb_data = 255;
12'd482 : rgb_data = 255;
12'd483 : rgb_data = 255;
12'd484 : rgb_data = 0;
12'd485 : rgb_data = 0;
12'd486 : rgb_data = 0;
12'd487 : rgb_data = 0;
12'd488 : rgb_data = 0;
12'd489 : rgb_data = 0;
12'd490 : rgb_data = 0;
12'd491 : rgb_data = 0;
12'd492 : rgb_data = 0;
12'd493 : rgb_data = 0;
12'd494 : rgb_data = 0;
12'd495 : rgb_data = 0;
12'd496 : rgb_data = 0;
12'd497 : rgb_data = 0;
12'd498 : rgb_data = 0;
12'd499 : rgb_data = 0;
12'd500 : rgb_data = 0;
12'd501 : rgb_data = 0;
12'd502 : rgb_data = 0;
12'd503 : rgb_data = 0;
12'd504 : rgb_data = 0;
12'd505 : rgb_data = 0;
12'd506 : rgb_data = 0;
12'd507 : rgb_data = 0;
12'd508 : rgb_data = 0;
12'd509 : rgb_data = 0;
12'd510 : rgb_data = 0;
12'd511 : rgb_data = 0;
12'd512 : rgb_data = 0;
12'd513 : rgb_data = 0;
12'd514 : rgb_data = 0;
12'd515 : rgb_data = 0;
12'd516 : rgb_data = 0;
12'd517 : rgb_data = 0;
12'd518 : rgb_data = 0;
12'd519 : rgb_data = 0;
12'd520 : rgb_data = 0;
12'd521 : rgb_data = 0;
12'd522 : rgb_data = 0;
12'd523 : rgb_data = 0;
12'd524 : rgb_data = 0;
12'd525 : rgb_data = 0;
12'd526 : rgb_data = 0;
12'd527 : rgb_data = 0;
12'd528 : rgb_data = 0;
12'd529 : rgb_data = 0;
12'd530 : rgb_data = 0;
12'd531 : rgb_data = 0;
12'd532 : rgb_data = 0;
12'd533 : rgb_data = 0;
12'd534 : rgb_data = 0;
12'd535 : rgb_data = 0;
12'd536 : rgb_data = 0;
12'd537 : rgb_data = 0;
12'd538 : rgb_data = 0;
12'd539 : rgb_data = 0;
12'd540 : rgb_data = 255;
12'd541 : rgb_data = 255;
12'd542 : rgb_data = 255;
12'd543 : rgb_data = 255;
12'd544 : rgb_data = 255;
12'd545 : rgb_data = 255;
12'd546 : rgb_data = 255;
12'd547 : rgb_data = 255;
12'd548 : rgb_data = 0;
12'd549 : rgb_data = 0;
12'd550 : rgb_data = 0;
12'd551 : rgb_data = 0;
12'd552 : rgb_data = 0;
12'd553 : rgb_data = 0;
12'd554 : rgb_data = 0;
12'd555 : rgb_data = 0;
12'd556 : rgb_data = 0;
12'd557 : rgb_data = 0;
12'd558 : rgb_data = 0;
12'd559 : rgb_data = 0;
12'd560 : rgb_data = 0;
12'd561 : rgb_data = 0;
12'd562 : rgb_data = 0;
12'd563 : rgb_data = 0;
12'd564 : rgb_data = 0;
12'd565 : rgb_data = 0;
12'd566 : rgb_data = 0;
12'd567 : rgb_data = 0;
12'd568 : rgb_data = 0;
12'd569 : rgb_data = 0;
12'd570 : rgb_data = 0;
12'd571 : rgb_data = 0;
12'd572 : rgb_data = 0;
12'd573 : rgb_data = 0;
12'd574 : rgb_data = 0;
12'd575 : rgb_data = 0;
12'd576 : rgb_data = 0;
12'd577 : rgb_data = 0;
12'd578 : rgb_data = 0;
12'd579 : rgb_data = 0;
12'd580 : rgb_data = 0;
12'd581 : rgb_data = 0;
12'd582 : rgb_data = 0;
12'd583 : rgb_data = 0;
12'd584 : rgb_data = 0;
12'd585 : rgb_data = 0;
12'd586 : rgb_data = 0;
12'd587 : rgb_data = 0;
12'd588 : rgb_data = 0;
12'd589 : rgb_data = 0;
12'd590 : rgb_data = 0;
12'd591 : rgb_data = 0;
12'd592 : rgb_data = 0;
12'd593 : rgb_data = 0;
12'd594 : rgb_data = 0;
12'd595 : rgb_data = 0;
12'd596 : rgb_data = 0;
12'd597 : rgb_data = 0;
12'd598 : rgb_data = 0;
12'd599 : rgb_data = 0;
12'd600 : rgb_data = 0;
12'd601 : rgb_data = 0;
12'd602 : rgb_data = 0;
12'd603 : rgb_data = 0;
12'd604 : rgb_data = 255;
12'd605 : rgb_data = 255;
12'd606 : rgb_data = 255;
12'd607 : rgb_data = 255;
12'd608 : rgb_data = 255;
12'd609 : rgb_data = 255;
12'd610 : rgb_data = 255;
12'd611 : rgb_data = 255;
12'd612 : rgb_data = 0;
12'd613 : rgb_data = 0;
12'd614 : rgb_data = 0;
12'd615 : rgb_data = 0;
12'd616 : rgb_data = 0;
12'd617 : rgb_data = 0;
12'd618 : rgb_data = 0;
12'd619 : rgb_data = 0;
12'd620 : rgb_data = 0;
12'd621 : rgb_data = 0;
12'd622 : rgb_data = 0;
12'd623 : rgb_data = 0;
12'd624 : rgb_data = 0;
12'd625 : rgb_data = 0;
12'd626 : rgb_data = 0;
12'd627 : rgb_data = 0;
12'd628 : rgb_data = 0;
12'd629 : rgb_data = 0;
12'd630 : rgb_data = 0;
12'd631 : rgb_data = 0;
12'd632 : rgb_data = 0;
12'd633 : rgb_data = 0;
12'd634 : rgb_data = 0;
12'd635 : rgb_data = 0;
12'd636 : rgb_data = 0;
12'd637 : rgb_data = 0;
12'd638 : rgb_data = 0;
12'd639 : rgb_data = 0;
12'd640 : rgb_data = 0;
12'd641 : rgb_data = 0;
12'd642 : rgb_data = 0;
12'd643 : rgb_data = 0;
12'd644 : rgb_data = 0;
12'd645 : rgb_data = 0;
12'd646 : rgb_data = 0;
12'd647 : rgb_data = 0;
12'd648 : rgb_data = 0;
12'd649 : rgb_data = 0;
12'd650 : rgb_data = 0;
12'd651 : rgb_data = 0;
12'd652 : rgb_data = 0;
12'd653 : rgb_data = 0;
12'd654 : rgb_data = 0;
12'd655 : rgb_data = 0;
12'd656 : rgb_data = 0;
12'd657 : rgb_data = 0;
12'd658 : rgb_data = 0;
12'd659 : rgb_data = 0;
12'd660 : rgb_data = 0;
12'd661 : rgb_data = 0;
12'd662 : rgb_data = 0;
12'd663 : rgb_data = 0;
12'd664 : rgb_data = 0;
12'd665 : rgb_data = 0;
12'd666 : rgb_data = 0;
12'd667 : rgb_data = 0;
12'd668 : rgb_data = 255;
12'd669 : rgb_data = 255;
12'd670 : rgb_data = 255;
12'd671 : rgb_data = 255;
12'd672 : rgb_data = 255;
12'd673 : rgb_data = 255;
12'd674 : rgb_data = 255;
12'd675 : rgb_data = 255;
12'd676 : rgb_data = 0;
12'd677 : rgb_data = 0;
12'd678 : rgb_data = 0;
12'd679 : rgb_data = 0;
12'd680 : rgb_data = 0;
12'd681 : rgb_data = 0;
12'd682 : rgb_data = 0;
12'd683 : rgb_data = 0;
12'd684 : rgb_data = 0;
12'd685 : rgb_data = 0;
12'd686 : rgb_data = 0;
12'd687 : rgb_data = 0;
12'd688 : rgb_data = 0;
12'd689 : rgb_data = 0;
12'd690 : rgb_data = 0;
12'd691 : rgb_data = 0;
12'd692 : rgb_data = 0;
12'd693 : rgb_data = 0;
12'd694 : rgb_data = 0;
12'd695 : rgb_data = 0;
12'd696 : rgb_data = 0;
12'd697 : rgb_data = 0;
12'd698 : rgb_data = 0;
12'd699 : rgb_data = 0;
12'd700 : rgb_data = 0;
12'd701 : rgb_data = 0;
12'd702 : rgb_data = 0;
12'd703 : rgb_data = 0;
12'd704 : rgb_data = 0;
12'd705 : rgb_data = 0;
12'd706 : rgb_data = 0;
12'd707 : rgb_data = 0;
12'd708 : rgb_data = 0;
12'd709 : rgb_data = 0;
12'd710 : rgb_data = 0;
12'd711 : rgb_data = 0;
12'd712 : rgb_data = 0;
12'd713 : rgb_data = 0;
12'd714 : rgb_data = 0;
12'd715 : rgb_data = 0;
12'd716 : rgb_data = 0;
12'd717 : rgb_data = 0;
12'd718 : rgb_data = 0;
12'd719 : rgb_data = 0;
12'd720 : rgb_data = 0;
12'd721 : rgb_data = 0;
12'd722 : rgb_data = 0;
12'd723 : rgb_data = 0;
12'd724 : rgb_data = 0;
12'd725 : rgb_data = 0;
12'd726 : rgb_data = 0;
12'd727 : rgb_data = 0;
12'd728 : rgb_data = 0;
12'd729 : rgb_data = 0;
12'd730 : rgb_data = 0;
12'd731 : rgb_data = 0;
12'd732 : rgb_data = 255;
12'd733 : rgb_data = 255;
12'd734 : rgb_data = 255;
12'd735 : rgb_data = 255;
12'd736 : rgb_data = 255;
12'd737 : rgb_data = 255;
12'd738 : rgb_data = 255;
12'd739 : rgb_data = 255;
12'd740 : rgb_data = 0;
12'd741 : rgb_data = 0;
12'd742 : rgb_data = 0;
12'd743 : rgb_data = 0;
12'd744 : rgb_data = 0;
12'd745 : rgb_data = 0;
12'd746 : rgb_data = 0;
12'd747 : rgb_data = 0;
12'd748 : rgb_data = 0;
12'd749 : rgb_data = 0;
12'd750 : rgb_data = 0;
12'd751 : rgb_data = 0;
12'd752 : rgb_data = 0;
12'd753 : rgb_data = 0;
12'd754 : rgb_data = 0;
12'd755 : rgb_data = 0;
12'd756 : rgb_data = 0;
12'd757 : rgb_data = 0;
12'd758 : rgb_data = 0;
12'd759 : rgb_data = 0;
12'd760 : rgb_data = 0;
12'd761 : rgb_data = 0;
12'd762 : rgb_data = 0;
12'd763 : rgb_data = 0;
12'd764 : rgb_data = 0;
12'd765 : rgb_data = 0;
12'd766 : rgb_data = 0;
12'd767 : rgb_data = 0;
12'd768 : rgb_data = 0;
12'd769 : rgb_data = 0;
12'd770 : rgb_data = 0;
12'd771 : rgb_data = 0;
12'd772 : rgb_data = 0;
12'd773 : rgb_data = 0;
12'd774 : rgb_data = 0;
12'd775 : rgb_data = 0;
12'd776 : rgb_data = 0;
12'd777 : rgb_data = 0;
12'd778 : rgb_data = 0;
12'd779 : rgb_data = 0;
12'd780 : rgb_data = 0;
12'd781 : rgb_data = 0;
12'd782 : rgb_data = 0;
12'd783 : rgb_data = 0;
12'd784 : rgb_data = 0;
12'd785 : rgb_data = 0;
12'd786 : rgb_data = 0;
12'd787 : rgb_data = 0;
12'd788 : rgb_data = 0;
12'd789 : rgb_data = 0;
12'd790 : rgb_data = 0;
12'd791 : rgb_data = 0;
12'd792 : rgb_data = 0;
12'd793 : rgb_data = 0;
12'd794 : rgb_data = 0;
12'd795 : rgb_data = 0;
12'd796 : rgb_data = 255;
12'd797 : rgb_data = 255;
12'd798 : rgb_data = 255;
12'd799 : rgb_data = 255;
12'd800 : rgb_data = 255;
12'd801 : rgb_data = 255;
12'd802 : rgb_data = 255;
12'd803 : rgb_data = 255;
12'd804 : rgb_data = 0;
12'd805 : rgb_data = 0;
12'd806 : rgb_data = 0;
12'd807 : rgb_data = 0;
12'd808 : rgb_data = 0;
12'd809 : rgb_data = 0;
12'd810 : rgb_data = 0;
12'd811 : rgb_data = 0;
12'd812 : rgb_data = 0;
12'd813 : rgb_data = 0;
12'd814 : rgb_data = 0;
12'd815 : rgb_data = 0;
12'd816 : rgb_data = 0;
12'd817 : rgb_data = 0;
12'd818 : rgb_data = 0;
12'd819 : rgb_data = 0;
12'd820 : rgb_data = 0;
12'd821 : rgb_data = 0;
12'd822 : rgb_data = 0;
12'd823 : rgb_data = 0;
12'd824 : rgb_data = 0;
12'd825 : rgb_data = 0;
12'd826 : rgb_data = 0;
12'd827 : rgb_data = 0;
12'd828 : rgb_data = 0;
12'd829 : rgb_data = 0;
12'd830 : rgb_data = 0;
12'd831 : rgb_data = 0;
12'd832 : rgb_data = 0;
12'd833 : rgb_data = 0;
12'd834 : rgb_data = 0;
12'd835 : rgb_data = 0;
12'd836 : rgb_data = 0;
12'd837 : rgb_data = 0;
12'd838 : rgb_data = 0;
12'd839 : rgb_data = 0;
12'd840 : rgb_data = 0;
12'd841 : rgb_data = 0;
12'd842 : rgb_data = 0;
12'd843 : rgb_data = 0;
12'd844 : rgb_data = 0;
12'd845 : rgb_data = 0;
12'd846 : rgb_data = 0;
12'd847 : rgb_data = 0;
12'd848 : rgb_data = 0;
12'd849 : rgb_data = 0;
12'd850 : rgb_data = 0;
12'd851 : rgb_data = 0;
12'd852 : rgb_data = 0;
12'd853 : rgb_data = 0;
12'd854 : rgb_data = 0;
12'd855 : rgb_data = 0;
12'd856 : rgb_data = 0;
12'd857 : rgb_data = 0;
12'd858 : rgb_data = 0;
12'd859 : rgb_data = 0;
12'd860 : rgb_data = 255;
12'd861 : rgb_data = 255;
12'd862 : rgb_data = 255;
12'd863 : rgb_data = 255;
12'd864 : rgb_data = 255;
12'd865 : rgb_data = 255;
12'd866 : rgb_data = 255;
12'd867 : rgb_data = 255;
12'd868 : rgb_data = 0;
12'd869 : rgb_data = 0;
12'd870 : rgb_data = 0;
12'd871 : rgb_data = 0;
12'd872 : rgb_data = 0;
12'd873 : rgb_data = 0;
12'd874 : rgb_data = 0;
12'd875 : rgb_data = 0;
12'd876 : rgb_data = 0;
12'd877 : rgb_data = 0;
12'd878 : rgb_data = 0;
12'd879 : rgb_data = 0;
12'd880 : rgb_data = 0;
12'd881 : rgb_data = 0;
12'd882 : rgb_data = 0;
12'd883 : rgb_data = 0;
12'd884 : rgb_data = 0;
12'd885 : rgb_data = 0;
12'd886 : rgb_data = 0;
12'd887 : rgb_data = 0;
12'd888 : rgb_data = 0;
12'd889 : rgb_data = 0;
12'd890 : rgb_data = 0;
12'd891 : rgb_data = 0;
12'd892 : rgb_data = 0;
12'd893 : rgb_data = 0;
12'd894 : rgb_data = 0;
12'd895 : rgb_data = 0;
12'd896 : rgb_data = 0;
12'd897 : rgb_data = 0;
12'd898 : rgb_data = 0;
12'd899 : rgb_data = 0;
12'd900 : rgb_data = 0;
12'd901 : rgb_data = 0;
12'd902 : rgb_data = 0;
12'd903 : rgb_data = 0;
12'd904 : rgb_data = 0;
12'd905 : rgb_data = 0;
12'd906 : rgb_data = 0;
12'd907 : rgb_data = 0;
12'd908 : rgb_data = 0;
12'd909 : rgb_data = 0;
12'd910 : rgb_data = 0;
12'd911 : rgb_data = 0;
12'd912 : rgb_data = 0;
12'd913 : rgb_data = 0;
12'd914 : rgb_data = 0;
12'd915 : rgb_data = 0;
12'd916 : rgb_data = 0;
12'd917 : rgb_data = 0;
12'd918 : rgb_data = 0;
12'd919 : rgb_data = 0;
12'd920 : rgb_data = 0;
12'd921 : rgb_data = 0;
12'd922 : rgb_data = 0;
12'd923 : rgb_data = 0;
12'd924 : rgb_data = 255;
12'd925 : rgb_data = 255;
12'd926 : rgb_data = 255;
12'd927 : rgb_data = 255;
12'd928 : rgb_data = 255;
12'd929 : rgb_data = 255;
12'd930 : rgb_data = 255;
12'd931 : rgb_data = 255;
12'd932 : rgb_data = 0;
12'd933 : rgb_data = 0;
12'd934 : rgb_data = 0;
12'd935 : rgb_data = 0;
12'd936 : rgb_data = 0;
12'd937 : rgb_data = 0;
12'd938 : rgb_data = 0;
12'd939 : rgb_data = 0;
12'd940 : rgb_data = 0;
12'd941 : rgb_data = 0;
12'd942 : rgb_data = 0;
12'd943 : rgb_data = 0;
12'd944 : rgb_data = 0;
12'd945 : rgb_data = 0;
12'd946 : rgb_data = 0;
12'd947 : rgb_data = 0;
12'd948 : rgb_data = 0;
12'd949 : rgb_data = 0;
12'd950 : rgb_data = 0;
12'd951 : rgb_data = 0;
12'd952 : rgb_data = 0;
12'd953 : rgb_data = 0;
12'd954 : rgb_data = 0;
12'd955 : rgb_data = 0;
12'd956 : rgb_data = 0;
12'd957 : rgb_data = 0;
12'd958 : rgb_data = 0;
12'd959 : rgb_data = 0;
12'd960 : rgb_data = 0;
12'd961 : rgb_data = 0;
12'd962 : rgb_data = 0;
12'd963 : rgb_data = 0;
12'd964 : rgb_data = 0;
12'd965 : rgb_data = 0;
12'd966 : rgb_data = 0;
12'd967 : rgb_data = 0;
12'd968 : rgb_data = 0;
12'd969 : rgb_data = 0;
12'd970 : rgb_data = 0;
12'd971 : rgb_data = 0;
12'd972 : rgb_data = 0;
12'd973 : rgb_data = 0;
12'd974 : rgb_data = 0;
12'd975 : rgb_data = 0;
12'd976 : rgb_data = 0;
12'd977 : rgb_data = 0;
12'd978 : rgb_data = 0;
12'd979 : rgb_data = 0;
12'd980 : rgb_data = 0;
12'd981 : rgb_data = 0;
12'd982 : rgb_data = 0;
12'd983 : rgb_data = 0;
12'd984 : rgb_data = 0;
12'd985 : rgb_data = 0;
12'd986 : rgb_data = 0;
12'd987 : rgb_data = 0;
12'd988 : rgb_data = 255;
12'd989 : rgb_data = 255;
12'd990 : rgb_data = 255;
12'd991 : rgb_data = 255;
12'd992 : rgb_data = 255;
12'd993 : rgb_data = 255;
12'd994 : rgb_data = 255;
12'd995 : rgb_data = 255;
12'd996 : rgb_data = 0;
12'd997 : rgb_data = 0;
12'd998 : rgb_data = 0;
12'd999 : rgb_data = 0;
12'd1000: rgb_data = 0;
12'd1001: rgb_data = 0;
12'd1002: rgb_data = 0;
12'd1003: rgb_data = 0;
12'd1004: rgb_data = 0;
12'd1005: rgb_data = 0;
12'd1006: rgb_data = 0;
12'd1007: rgb_data = 0;
12'd1008: rgb_data = 0;
12'd1009: rgb_data = 0;
12'd1010: rgb_data = 0;
12'd1011: rgb_data = 0;
12'd1012: rgb_data = 0;
12'd1013: rgb_data = 0;
12'd1014: rgb_data = 0;
12'd1015: rgb_data = 0;
12'd1016: rgb_data = 0;
12'd1017: rgb_data = 0;
12'd1018: rgb_data = 0;
12'd1019: rgb_data = 0;
12'd1020: rgb_data = 0;
12'd1021: rgb_data = 0;
12'd1022: rgb_data = 0;
12'd1023: rgb_data = 0;
12'd1024: rgb_data = 0;
12'd1025: rgb_data = 0;
12'd1026: rgb_data = 0;
12'd1027: rgb_data = 0;
12'd1028: rgb_data = 0;
12'd1029: rgb_data = 0;
12'd1030: rgb_data = 0;
12'd1031: rgb_data = 0;
12'd1032: rgb_data = 0;
12'd1033: rgb_data = 0;
12'd1034: rgb_data = 0;
12'd1035: rgb_data = 0;
12'd1036: rgb_data = 0;
12'd1037: rgb_data = 0;
12'd1038: rgb_data = 0;
12'd1039: rgb_data = 0;
12'd1040: rgb_data = 0;
12'd1041: rgb_data = 0;
12'd1042: rgb_data = 0;
12'd1043: rgb_data = 0;
12'd1044: rgb_data = 0;
12'd1045: rgb_data = 0;
12'd1046: rgb_data = 0;
12'd1047: rgb_data = 0;
12'd1048: rgb_data = 0;
12'd1049: rgb_data = 0;
12'd1050: rgb_data = 0;
12'd1051: rgb_data = 0;
12'd1052: rgb_data = 255;
12'd1053: rgb_data = 255;
12'd1054: rgb_data = 255;
12'd1055: rgb_data = 255;
12'd1056: rgb_data = 255;
12'd1057: rgb_data = 255;
12'd1058: rgb_data = 255;
12'd1059: rgb_data = 255;
12'd1060: rgb_data = 0;
12'd1061: rgb_data = 0;
12'd1062: rgb_data = 0;
12'd1063: rgb_data = 0;
12'd1064: rgb_data = 0;
12'd1065: rgb_data = 0;
12'd1066: rgb_data = 0;
12'd1067: rgb_data = 0;
12'd1068: rgb_data = 0;
12'd1069: rgb_data = 0;
12'd1070: rgb_data = 0;
12'd1071: rgb_data = 0;
12'd1072: rgb_data = 0;
12'd1073: rgb_data = 0;
12'd1074: rgb_data = 0;
12'd1075: rgb_data = 0;
12'd1076: rgb_data = 0;
12'd1077: rgb_data = 0;
12'd1078: rgb_data = 0;
12'd1079: rgb_data = 0;
12'd1080: rgb_data = 0;
12'd1081: rgb_data = 0;
12'd1082: rgb_data = 0;
12'd1083: rgb_data = 0;
12'd1084: rgb_data = 0;
12'd1085: rgb_data = 0;
12'd1086: rgb_data = 0;
12'd1087: rgb_data = 0;
12'd1088: rgb_data = 0;
12'd1089: rgb_data = 0;
12'd1090: rgb_data = 0;
12'd1091: rgb_data = 0;
12'd1092: rgb_data = 0;
12'd1093: rgb_data = 0;
12'd1094: rgb_data = 0;
12'd1095: rgb_data = 0;
12'd1096: rgb_data = 0;
12'd1097: rgb_data = 0;
12'd1098: rgb_data = 0;
12'd1099: rgb_data = 0;
12'd1100: rgb_data = 0;
12'd1101: rgb_data = 0;
12'd1102: rgb_data = 0;
12'd1103: rgb_data = 0;
12'd1104: rgb_data = 0;
12'd1105: rgb_data = 0;
12'd1106: rgb_data = 0;
12'd1107: rgb_data = 0;
12'd1108: rgb_data = 0;
12'd1109: rgb_data = 0;
12'd1110: rgb_data = 0;
12'd1111: rgb_data = 0;
12'd1112: rgb_data = 0;
12'd1113: rgb_data = 0;
12'd1114: rgb_data = 0;
12'd1115: rgb_data = 0;
12'd1116: rgb_data = 255;
12'd1117: rgb_data = 255;
12'd1118: rgb_data = 255;
12'd1119: rgb_data = 255;
12'd1120: rgb_data = 255;
12'd1121: rgb_data = 255;
12'd1122: rgb_data = 255;
12'd1123: rgb_data = 255;
12'd1124: rgb_data = 0;
12'd1125: rgb_data = 0;
12'd1126: rgb_data = 0;
12'd1127: rgb_data = 0;
12'd1128: rgb_data = 0;
12'd1129: rgb_data = 0;
12'd1130: rgb_data = 0;
12'd1131: rgb_data = 0;
12'd1132: rgb_data = 0;
12'd1133: rgb_data = 0;
12'd1134: rgb_data = 0;
12'd1135: rgb_data = 0;
12'd1136: rgb_data = 0;
12'd1137: rgb_data = 0;
12'd1138: rgb_data = 0;
12'd1139: rgb_data = 0;
12'd1140: rgb_data = 0;
12'd1141: rgb_data = 0;
12'd1142: rgb_data = 0;
12'd1143: rgb_data = 0;
12'd1144: rgb_data = 0;
12'd1145: rgb_data = 0;
12'd1146: rgb_data = 0;
12'd1147: rgb_data = 0;
12'd1148: rgb_data = 0;
12'd1149: rgb_data = 0;
12'd1150: rgb_data = 0;
12'd1151: rgb_data = 0;
12'd1152: rgb_data = 0;
12'd1153: rgb_data = 0;
12'd1154: rgb_data = 0;
12'd1155: rgb_data = 0;
12'd1156: rgb_data = 0;
12'd1157: rgb_data = 0;
12'd1158: rgb_data = 0;
12'd1159: rgb_data = 0;
12'd1160: rgb_data = 0;
12'd1161: rgb_data = 0;
12'd1162: rgb_data = 0;
12'd1163: rgb_data = 0;
12'd1164: rgb_data = 0;
12'd1165: rgb_data = 0;
12'd1166: rgb_data = 0;
12'd1167: rgb_data = 0;
12'd1168: rgb_data = 0;
12'd1169: rgb_data = 0;
12'd1170: rgb_data = 0;
12'd1171: rgb_data = 0;
12'd1172: rgb_data = 0;
12'd1173: rgb_data = 0;
12'd1174: rgb_data = 0;
12'd1175: rgb_data = 0;
12'd1176: rgb_data = 0;
12'd1177: rgb_data = 0;
12'd1178: rgb_data = 0;
12'd1179: rgb_data = 0;
12'd1180: rgb_data = 255;
12'd1181: rgb_data = 255;
12'd1182: rgb_data = 255;
12'd1183: rgb_data = 255;
12'd1184: rgb_data = 255;
12'd1185: rgb_data = 255;
12'd1186: rgb_data = 255;
12'd1187: rgb_data = 255;
12'd1188: rgb_data = 0;
12'd1189: rgb_data = 0;
12'd1190: rgb_data = 0;
12'd1191: rgb_data = 0;
12'd1192: rgb_data = 0;
12'd1193: rgb_data = 0;
12'd1194: rgb_data = 0;
12'd1195: rgb_data = 0;
12'd1196: rgb_data = 0;
12'd1197: rgb_data = 0;
12'd1198: rgb_data = 0;
12'd1199: rgb_data = 0;
12'd1200: rgb_data = 0;
12'd1201: rgb_data = 0;
12'd1202: rgb_data = 0;
12'd1203: rgb_data = 0;
12'd1204: rgb_data = 0;
12'd1205: rgb_data = 0;
12'd1206: rgb_data = 0;
12'd1207: rgb_data = 0;
12'd1208: rgb_data = 0;
12'd1209: rgb_data = 0;
12'd1210: rgb_data = 0;
12'd1211: rgb_data = 0;
12'd1212: rgb_data = 0;
12'd1213: rgb_data = 0;
12'd1214: rgb_data = 0;
12'd1215: rgb_data = 0;
12'd1216: rgb_data = 0;
12'd1217: rgb_data = 0;
12'd1218: rgb_data = 0;
12'd1219: rgb_data = 0;
12'd1220: rgb_data = 0;
12'd1221: rgb_data = 0;
12'd1222: rgb_data = 0;
12'd1223: rgb_data = 0;
12'd1224: rgb_data = 0;
12'd1225: rgb_data = 0;
12'd1226: rgb_data = 0;
12'd1227: rgb_data = 0;
12'd1228: rgb_data = 0;
12'd1229: rgb_data = 0;
12'd1230: rgb_data = 0;
12'd1231: rgb_data = 0;
12'd1232: rgb_data = 0;
12'd1233: rgb_data = 0;
12'd1234: rgb_data = 0;
12'd1235: rgb_data = 0;
12'd1236: rgb_data = 0;
12'd1237: rgb_data = 0;
12'd1238: rgb_data = 0;
12'd1239: rgb_data = 0;
12'd1240: rgb_data = 0;
12'd1241: rgb_data = 0;
12'd1242: rgb_data = 0;
12'd1243: rgb_data = 0;
12'd1244: rgb_data = 255;
12'd1245: rgb_data = 255;
12'd1246: rgb_data = 255;
12'd1247: rgb_data = 255;
12'd1248: rgb_data = 255;
12'd1249: rgb_data = 255;
12'd1250: rgb_data = 255;
12'd1251: rgb_data = 255;
12'd1252: rgb_data = 0;
12'd1253: rgb_data = 0;
12'd1254: rgb_data = 0;
12'd1255: rgb_data = 0;
12'd1256: rgb_data = 0;
12'd1257: rgb_data = 0;
12'd1258: rgb_data = 0;
12'd1259: rgb_data = 0;
12'd1260: rgb_data = 0;
12'd1261: rgb_data = 0;
12'd1262: rgb_data = 0;
12'd1263: rgb_data = 0;
12'd1264: rgb_data = 0;
12'd1265: rgb_data = 0;
12'd1266: rgb_data = 0;
12'd1267: rgb_data = 0;
12'd1268: rgb_data = 0;
12'd1269: rgb_data = 0;
12'd1270: rgb_data = 0;
12'd1271: rgb_data = 0;
12'd1272: rgb_data = 0;
12'd1273: rgb_data = 0;
12'd1274: rgb_data = 0;
12'd1275: rgb_data = 0;
12'd1276: rgb_data = 0;
12'd1277: rgb_data = 0;
12'd1278: rgb_data = 0;
12'd1279: rgb_data = 0;
12'd1280: rgb_data = 0;
12'd1281: rgb_data = 0;
12'd1282: rgb_data = 0;
12'd1283: rgb_data = 0;
12'd1284: rgb_data = 0;
12'd1285: rgb_data = 0;
12'd1286: rgb_data = 0;
12'd1287: rgb_data = 0;
12'd1288: rgb_data = 0;
12'd1289: rgb_data = 0;
12'd1290: rgb_data = 0;
12'd1291: rgb_data = 0;
12'd1292: rgb_data = 0;
12'd1293: rgb_data = 0;
12'd1294: rgb_data = 0;
12'd1295: rgb_data = 0;
12'd1296: rgb_data = 0;
12'd1297: rgb_data = 0;
12'd1298: rgb_data = 0;
12'd1299: rgb_data = 0;
12'd1300: rgb_data = 0;
12'd1301: rgb_data = 0;
12'd1302: rgb_data = 0;
12'd1303: rgb_data = 0;
12'd1304: rgb_data = 0;
12'd1305: rgb_data = 0;
12'd1306: rgb_data = 0;
12'd1307: rgb_data = 0;
12'd1308: rgb_data = 255;
12'd1309: rgb_data = 255;
12'd1310: rgb_data = 255;
12'd1311: rgb_data = 255;
12'd1312: rgb_data = 255;
12'd1313: rgb_data = 255;
12'd1314: rgb_data = 255;
12'd1315: rgb_data = 255;
12'd1316: rgb_data = 0;
12'd1317: rgb_data = 0;
12'd1318: rgb_data = 0;
12'd1319: rgb_data = 0;
12'd1320: rgb_data = 0;
12'd1321: rgb_data = 0;
12'd1322: rgb_data = 0;
12'd1323: rgb_data = 0;
12'd1324: rgb_data = 0;
12'd1325: rgb_data = 0;
12'd1326: rgb_data = 0;
12'd1327: rgb_data = 0;
12'd1328: rgb_data = 0;
12'd1329: rgb_data = 0;
12'd1330: rgb_data = 0;
12'd1331: rgb_data = 0;
12'd1332: rgb_data = 0;
12'd1333: rgb_data = 0;
12'd1334: rgb_data = 0;
12'd1335: rgb_data = 0;
12'd1336: rgb_data = 0;
12'd1337: rgb_data = 0;
12'd1338: rgb_data = 0;
12'd1339: rgb_data = 0;
12'd1340: rgb_data = 0;
12'd1341: rgb_data = 0;
12'd1342: rgb_data = 0;
12'd1343: rgb_data = 0;
12'd1344: rgb_data = 0;
12'd1345: rgb_data = 0;
12'd1346: rgb_data = 0;
12'd1347: rgb_data = 0;
12'd1348: rgb_data = 0;
12'd1349: rgb_data = 0;
12'd1350: rgb_data = 0;
12'd1351: rgb_data = 0;
12'd1352: rgb_data = 0;
12'd1353: rgb_data = 0;
12'd1354: rgb_data = 0;
12'd1355: rgb_data = 0;
12'd1356: rgb_data = 0;
12'd1357: rgb_data = 0;
12'd1358: rgb_data = 0;
12'd1359: rgb_data = 0;
12'd1360: rgb_data = 0;
12'd1361: rgb_data = 0;
12'd1362: rgb_data = 0;
12'd1363: rgb_data = 0;
12'd1364: rgb_data = 0;
12'd1365: rgb_data = 0;
12'd1366: rgb_data = 0;
12'd1367: rgb_data = 0;
12'd1368: rgb_data = 0;
12'd1369: rgb_data = 0;
12'd1370: rgb_data = 0;
12'd1371: rgb_data = 0;
12'd1372: rgb_data = 255;
12'd1373: rgb_data = 255;
12'd1374: rgb_data = 255;
12'd1375: rgb_data = 255;
12'd1376: rgb_data = 255;
12'd1377: rgb_data = 255;
12'd1378: rgb_data = 255;
12'd1379: rgb_data = 255;
12'd1380: rgb_data = 0;
12'd1381: rgb_data = 0;
12'd1382: rgb_data = 0;
12'd1383: rgb_data = 0;
12'd1384: rgb_data = 0;
12'd1385: rgb_data = 0;
12'd1386: rgb_data = 0;
12'd1387: rgb_data = 0;
12'd1388: rgb_data = 0;
12'd1389: rgb_data = 0;
12'd1390: rgb_data = 0;
12'd1391: rgb_data = 0;
12'd1392: rgb_data = 0;
12'd1393: rgb_data = 0;
12'd1394: rgb_data = 0;
12'd1395: rgb_data = 0;
12'd1396: rgb_data = 0;
12'd1397: rgb_data = 0;
12'd1398: rgb_data = 0;
12'd1399: rgb_data = 0;
12'd1400: rgb_data = 0;
12'd1401: rgb_data = 0;
12'd1402: rgb_data = 0;
12'd1403: rgb_data = 0;
12'd1404: rgb_data = 0;
12'd1405: rgb_data = 0;
12'd1406: rgb_data = 0;
12'd1407: rgb_data = 0;
12'd1408: rgb_data = 0;
12'd1409: rgb_data = 0;
12'd1410: rgb_data = 0;
12'd1411: rgb_data = 0;
12'd1412: rgb_data = 0;
12'd1413: rgb_data = 0;
12'd1414: rgb_data = 0;
12'd1415: rgb_data = 0;
12'd1416: rgb_data = 0;
12'd1417: rgb_data = 0;
12'd1418: rgb_data = 0;
12'd1419: rgb_data = 0;
12'd1420: rgb_data = 0;
12'd1421: rgb_data = 0;
12'd1422: rgb_data = 0;
12'd1423: rgb_data = 0;
12'd1424: rgb_data = 0;
12'd1425: rgb_data = 0;
12'd1426: rgb_data = 0;
12'd1427: rgb_data = 0;
12'd1428: rgb_data = 0;
12'd1429: rgb_data = 0;
12'd1430: rgb_data = 0;
12'd1431: rgb_data = 0;
12'd1432: rgb_data = 0;
12'd1433: rgb_data = 0;
12'd1434: rgb_data = 0;
12'd1435: rgb_data = 0;
12'd1436: rgb_data = 255;
12'd1437: rgb_data = 255;
12'd1438: rgb_data = 255;
12'd1439: rgb_data = 255;
12'd1440: rgb_data = 255;
12'd1441: rgb_data = 255;
12'd1442: rgb_data = 255;
12'd1443: rgb_data = 255;
12'd1444: rgb_data = 0;
12'd1445: rgb_data = 0;
12'd1446: rgb_data = 0;
12'd1447: rgb_data = 0;
12'd1448: rgb_data = 0;
12'd1449: rgb_data = 0;
12'd1450: rgb_data = 0;
12'd1451: rgb_data = 0;
12'd1452: rgb_data = 0;
12'd1453: rgb_data = 0;
12'd1454: rgb_data = 0;
12'd1455: rgb_data = 0;
12'd1456: rgb_data = 0;
12'd1457: rgb_data = 0;
12'd1458: rgb_data = 0;
12'd1459: rgb_data = 0;
12'd1460: rgb_data = 0;
12'd1461: rgb_data = 0;
12'd1462: rgb_data = 0;
12'd1463: rgb_data = 0;
12'd1464: rgb_data = 0;
12'd1465: rgb_data = 0;
12'd1466: rgb_data = 0;
12'd1467: rgb_data = 0;
12'd1468: rgb_data = 0;
12'd1469: rgb_data = 0;
12'd1470: rgb_data = 0;
12'd1471: rgb_data = 0;
12'd1472: rgb_data = 0;
12'd1473: rgb_data = 0;
12'd1474: rgb_data = 0;
12'd1475: rgb_data = 0;
12'd1476: rgb_data = 0;
12'd1477: rgb_data = 0;
12'd1478: rgb_data = 0;
12'd1479: rgb_data = 0;
12'd1480: rgb_data = 0;
12'd1481: rgb_data = 0;
12'd1482: rgb_data = 0;
12'd1483: rgb_data = 0;
12'd1484: rgb_data = 0;
12'd1485: rgb_data = 0;
12'd1486: rgb_data = 0;
12'd1487: rgb_data = 0;
12'd1488: rgb_data = 0;
12'd1489: rgb_data = 0;
12'd1490: rgb_data = 0;
12'd1491: rgb_data = 0;
12'd1492: rgb_data = 0;
12'd1493: rgb_data = 0;
12'd1494: rgb_data = 0;
12'd1495: rgb_data = 0;
12'd1496: rgb_data = 0;
12'd1497: rgb_data = 0;
12'd1498: rgb_data = 0;
12'd1499: rgb_data = 0;
12'd1500: rgb_data = 255;
12'd1501: rgb_data = 255;
12'd1502: rgb_data = 255;
12'd1503: rgb_data = 255;
12'd1504: rgb_data = 255;
12'd1505: rgb_data = 255;
12'd1506: rgb_data = 255;
12'd1507: rgb_data = 255;
12'd1508: rgb_data = 0;
12'd1509: rgb_data = 0;
12'd1510: rgb_data = 0;
12'd1511: rgb_data = 0;
12'd1512: rgb_data = 0;
12'd1513: rgb_data = 0;
12'd1514: rgb_data = 0;
12'd1515: rgb_data = 0;
12'd1516: rgb_data = 0;
12'd1517: rgb_data = 0;
12'd1518: rgb_data = 0;
12'd1519: rgb_data = 0;
12'd1520: rgb_data = 0;
12'd1521: rgb_data = 0;
12'd1522: rgb_data = 0;
12'd1523: rgb_data = 0;
12'd1524: rgb_data = 0;
12'd1525: rgb_data = 0;
12'd1526: rgb_data = 0;
12'd1527: rgb_data = 0;
12'd1528: rgb_data = 0;
12'd1529: rgb_data = 0;
12'd1530: rgb_data = 0;
12'd1531: rgb_data = 0;
12'd1532: rgb_data = 0;
12'd1533: rgb_data = 0;
12'd1534: rgb_data = 0;
12'd1535: rgb_data = 0;
12'd1536: rgb_data = 0;
12'd1537: rgb_data = 0;
12'd1538: rgb_data = 0;
12'd1539: rgb_data = 0;
12'd1540: rgb_data = 0;
12'd1541: rgb_data = 0;
12'd1542: rgb_data = 0;
12'd1543: rgb_data = 0;
12'd1544: rgb_data = 0;
12'd1545: rgb_data = 0;
12'd1546: rgb_data = 0;
12'd1547: rgb_data = 0;
12'd1548: rgb_data = 228;
12'd1549: rgb_data = 228;
12'd1550: rgb_data = 228;
12'd1551: rgb_data = 228;
12'd1552: rgb_data = 0;
12'd1553: rgb_data = 0;
12'd1554: rgb_data = 0;
12'd1555: rgb_data = 0;
12'd1556: rgb_data = 0;
12'd1557: rgb_data = 0;
12'd1558: rgb_data = 0;
12'd1559: rgb_data = 0;
12'd1560: rgb_data = 255;
12'd1561: rgb_data = 255;
12'd1562: rgb_data = 255;
12'd1563: rgb_data = 255;
12'd1564: rgb_data = 255;
12'd1565: rgb_data = 255;
12'd1566: rgb_data = 255;
12'd1567: rgb_data = 255;
12'd1568: rgb_data = 255;
12'd1569: rgb_data = 255;
12'd1570: rgb_data = 255;
12'd1571: rgb_data = 255;
12'd1572: rgb_data = 255;
12'd1573: rgb_data = 255;
12'd1574: rgb_data = 255;
12'd1575: rgb_data = 255;
12'd1576: rgb_data = 0;
12'd1577: rgb_data = 0;
12'd1578: rgb_data = 0;
12'd1579: rgb_data = 0;
12'd1580: rgb_data = 0;
12'd1581: rgb_data = 0;
12'd1582: rgb_data = 0;
12'd1583: rgb_data = 0;
12'd1584: rgb_data = 228;
12'd1585: rgb_data = 228;
12'd1586: rgb_data = 228;
12'd1587: rgb_data = 228;
12'd1588: rgb_data = 0;
12'd1589: rgb_data = 0;
12'd1590: rgb_data = 0;
12'd1591: rgb_data = 0;
12'd1592: rgb_data = 0;
12'd1593: rgb_data = 0;
12'd1594: rgb_data = 0;
12'd1595: rgb_data = 0;
12'd1596: rgb_data = 0;
12'd1597: rgb_data = 0;
12'd1598: rgb_data = 0;
12'd1599: rgb_data = 0;
12'd1600: rgb_data = 0;
12'd1601: rgb_data = 0;
12'd1602: rgb_data = 0;
12'd1603: rgb_data = 0;
12'd1604: rgb_data = 0;
12'd1605: rgb_data = 0;
12'd1606: rgb_data = 0;
12'd1607: rgb_data = 0;
12'd1608: rgb_data = 0;
12'd1609: rgb_data = 0;
12'd1610: rgb_data = 0;
12'd1611: rgb_data = 0;
12'd1612: rgb_data = 228;
12'd1613: rgb_data = 228;
12'd1614: rgb_data = 228;
12'd1615: rgb_data = 228;
12'd1616: rgb_data = 0;
12'd1617: rgb_data = 0;
12'd1618: rgb_data = 0;
12'd1619: rgb_data = 0;
12'd1620: rgb_data = 0;
12'd1621: rgb_data = 0;
12'd1622: rgb_data = 0;
12'd1623: rgb_data = 0;
12'd1624: rgb_data = 255;
12'd1625: rgb_data = 255;
12'd1626: rgb_data = 255;
12'd1627: rgb_data = 255;
12'd1628: rgb_data = 255;
12'd1629: rgb_data = 255;
12'd1630: rgb_data = 255;
12'd1631: rgb_data = 255;
12'd1632: rgb_data = 255;
12'd1633: rgb_data = 255;
12'd1634: rgb_data = 255;
12'd1635: rgb_data = 255;
12'd1636: rgb_data = 255;
12'd1637: rgb_data = 255;
12'd1638: rgb_data = 255;
12'd1639: rgb_data = 255;
12'd1640: rgb_data = 0;
12'd1641: rgb_data = 0;
12'd1642: rgb_data = 0;
12'd1643: rgb_data = 0;
12'd1644: rgb_data = 0;
12'd1645: rgb_data = 0;
12'd1646: rgb_data = 0;
12'd1647: rgb_data = 0;
12'd1648: rgb_data = 228;
12'd1649: rgb_data = 228;
12'd1650: rgb_data = 228;
12'd1651: rgb_data = 228;
12'd1652: rgb_data = 0;
12'd1653: rgb_data = 0;
12'd1654: rgb_data = 0;
12'd1655: rgb_data = 0;
12'd1656: rgb_data = 0;
12'd1657: rgb_data = 0;
12'd1658: rgb_data = 0;
12'd1659: rgb_data = 0;
12'd1660: rgb_data = 0;
12'd1661: rgb_data = 0;
12'd1662: rgb_data = 0;
12'd1663: rgb_data = 0;
12'd1664: rgb_data = 0;
12'd1665: rgb_data = 0;
12'd1666: rgb_data = 0;
12'd1667: rgb_data = 0;
12'd1668: rgb_data = 0;
12'd1669: rgb_data = 0;
12'd1670: rgb_data = 0;
12'd1671: rgb_data = 0;
12'd1672: rgb_data = 0;
12'd1673: rgb_data = 0;
12'd1674: rgb_data = 0;
12'd1675: rgb_data = 0;
12'd1676: rgb_data = 228;
12'd1677: rgb_data = 228;
12'd1678: rgb_data = 228;
12'd1679: rgb_data = 228;
12'd1680: rgb_data = 0;
12'd1681: rgb_data = 0;
12'd1682: rgb_data = 0;
12'd1683: rgb_data = 0;
12'd1684: rgb_data = 0;
12'd1685: rgb_data = 0;
12'd1686: rgb_data = 0;
12'd1687: rgb_data = 0;
12'd1688: rgb_data = 255;
12'd1689: rgb_data = 255;
12'd1690: rgb_data = 255;
12'd1691: rgb_data = 255;
12'd1692: rgb_data = 255;
12'd1693: rgb_data = 255;
12'd1694: rgb_data = 255;
12'd1695: rgb_data = 255;
12'd1696: rgb_data = 255;
12'd1697: rgb_data = 255;
12'd1698: rgb_data = 255;
12'd1699: rgb_data = 255;
12'd1700: rgb_data = 255;
12'd1701: rgb_data = 255;
12'd1702: rgb_data = 255;
12'd1703: rgb_data = 255;
12'd1704: rgb_data = 0;
12'd1705: rgb_data = 0;
12'd1706: rgb_data = 0;
12'd1707: rgb_data = 0;
12'd1708: rgb_data = 0;
12'd1709: rgb_data = 0;
12'd1710: rgb_data = 0;
12'd1711: rgb_data = 0;
12'd1712: rgb_data = 228;
12'd1713: rgb_data = 228;
12'd1714: rgb_data = 228;
12'd1715: rgb_data = 228;
12'd1716: rgb_data = 0;
12'd1717: rgb_data = 0;
12'd1718: rgb_data = 0;
12'd1719: rgb_data = 0;
12'd1720: rgb_data = 0;
12'd1721: rgb_data = 0;
12'd1722: rgb_data = 0;
12'd1723: rgb_data = 0;
12'd1724: rgb_data = 0;
12'd1725: rgb_data = 0;
12'd1726: rgb_data = 0;
12'd1727: rgb_data = 0;
12'd1728: rgb_data = 0;
12'd1729: rgb_data = 0;
12'd1730: rgb_data = 0;
12'd1731: rgb_data = 0;
12'd1732: rgb_data = 0;
12'd1733: rgb_data = 0;
12'd1734: rgb_data = 0;
12'd1735: rgb_data = 0;
12'd1736: rgb_data = 0;
12'd1737: rgb_data = 0;
12'd1738: rgb_data = 0;
12'd1739: rgb_data = 0;
12'd1740: rgb_data = 228;
12'd1741: rgb_data = 228;
12'd1742: rgb_data = 228;
12'd1743: rgb_data = 228;
12'd1744: rgb_data = 0;
12'd1745: rgb_data = 0;
12'd1746: rgb_data = 0;
12'd1747: rgb_data = 0;
12'd1748: rgb_data = 0;
12'd1749: rgb_data = 0;
12'd1750: rgb_data = 0;
12'd1751: rgb_data = 0;
12'd1752: rgb_data = 255;
12'd1753: rgb_data = 255;
12'd1754: rgb_data = 255;
12'd1755: rgb_data = 255;
12'd1756: rgb_data = 255;
12'd1757: rgb_data = 255;
12'd1758: rgb_data = 255;
12'd1759: rgb_data = 255;
12'd1760: rgb_data = 255;
12'd1761: rgb_data = 255;
12'd1762: rgb_data = 255;
12'd1763: rgb_data = 255;
12'd1764: rgb_data = 255;
12'd1765: rgb_data = 255;
12'd1766: rgb_data = 255;
12'd1767: rgb_data = 255;
12'd1768: rgb_data = 0;
12'd1769: rgb_data = 0;
12'd1770: rgb_data = 0;
12'd1771: rgb_data = 0;
12'd1772: rgb_data = 0;
12'd1773: rgb_data = 0;
12'd1774: rgb_data = 0;
12'd1775: rgb_data = 0;
12'd1776: rgb_data = 228;
12'd1777: rgb_data = 228;
12'd1778: rgb_data = 228;
12'd1779: rgb_data = 228;
12'd1780: rgb_data = 0;
12'd1781: rgb_data = 0;
12'd1782: rgb_data = 0;
12'd1783: rgb_data = 0;
12'd1784: rgb_data = 0;
12'd1785: rgb_data = 0;
12'd1786: rgb_data = 0;
12'd1787: rgb_data = 0;
12'd1788: rgb_data = 0;
12'd1789: rgb_data = 0;
12'd1790: rgb_data = 0;
12'd1791: rgb_data = 0;
12'd1792: rgb_data = 228;
12'd1793: rgb_data = 228;
12'd1794: rgb_data = 228;
12'd1795: rgb_data = 228;
12'd1796: rgb_data = 0;
12'd1797: rgb_data = 0;
12'd1798: rgb_data = 0;
12'd1799: rgb_data = 0;
12'd1800: rgb_data = 0;
12'd1801: rgb_data = 0;
12'd1802: rgb_data = 0;
12'd1803: rgb_data = 0;
12'd1804: rgb_data = 228;
12'd1805: rgb_data = 228;
12'd1806: rgb_data = 228;
12'd1807: rgb_data = 228;
12'd1808: rgb_data = 0;
12'd1809: rgb_data = 0;
12'd1810: rgb_data = 0;
12'd1811: rgb_data = 0;
12'd1812: rgb_data = 0;
12'd1813: rgb_data = 0;
12'd1814: rgb_data = 0;
12'd1815: rgb_data = 0;
12'd1816: rgb_data = 255;
12'd1817: rgb_data = 255;
12'd1818: rgb_data = 255;
12'd1819: rgb_data = 255;
12'd1820: rgb_data = 248;
12'd1821: rgb_data = 248;
12'd1822: rgb_data = 248;
12'd1823: rgb_data = 248;
12'd1824: rgb_data = 248;
12'd1825: rgb_data = 248;
12'd1826: rgb_data = 248;
12'd1827: rgb_data = 248;
12'd1828: rgb_data = 255;
12'd1829: rgb_data = 255;
12'd1830: rgb_data = 255;
12'd1831: rgb_data = 255;
12'd1832: rgb_data = 0;
12'd1833: rgb_data = 0;
12'd1834: rgb_data = 0;
12'd1835: rgb_data = 0;
12'd1836: rgb_data = 0;
12'd1837: rgb_data = 0;
12'd1838: rgb_data = 0;
12'd1839: rgb_data = 0;
12'd1840: rgb_data = 228;
12'd1841: rgb_data = 228;
12'd1842: rgb_data = 228;
12'd1843: rgb_data = 228;
12'd1844: rgb_data = 0;
12'd1845: rgb_data = 0;
12'd1846: rgb_data = 0;
12'd1847: rgb_data = 0;
12'd1848: rgb_data = 0;
12'd1849: rgb_data = 0;
12'd1850: rgb_data = 0;
12'd1851: rgb_data = 0;
12'd1852: rgb_data = 228;
12'd1853: rgb_data = 228;
12'd1854: rgb_data = 228;
12'd1855: rgb_data = 228;
12'd1856: rgb_data = 228;
12'd1857: rgb_data = 228;
12'd1858: rgb_data = 228;
12'd1859: rgb_data = 228;
12'd1860: rgb_data = 0;
12'd1861: rgb_data = 0;
12'd1862: rgb_data = 0;
12'd1863: rgb_data = 0;
12'd1864: rgb_data = 0;
12'd1865: rgb_data = 0;
12'd1866: rgb_data = 0;
12'd1867: rgb_data = 0;
12'd1868: rgb_data = 228;
12'd1869: rgb_data = 228;
12'd1870: rgb_data = 228;
12'd1871: rgb_data = 228;
12'd1872: rgb_data = 0;
12'd1873: rgb_data = 0;
12'd1874: rgb_data = 0;
12'd1875: rgb_data = 0;
12'd1876: rgb_data = 0;
12'd1877: rgb_data = 0;
12'd1878: rgb_data = 0;
12'd1879: rgb_data = 0;
12'd1880: rgb_data = 255;
12'd1881: rgb_data = 255;
12'd1882: rgb_data = 255;
12'd1883: rgb_data = 255;
12'd1884: rgb_data = 248;
12'd1885: rgb_data = 248;
12'd1886: rgb_data = 248;
12'd1887: rgb_data = 248;
12'd1888: rgb_data = 248;
12'd1889: rgb_data = 248;
12'd1890: rgb_data = 248;
12'd1891: rgb_data = 248;
12'd1892: rgb_data = 255;
12'd1893: rgb_data = 255;
12'd1894: rgb_data = 255;
12'd1895: rgb_data = 255;
12'd1896: rgb_data = 0;
12'd1897: rgb_data = 0;
12'd1898: rgb_data = 0;
12'd1899: rgb_data = 0;
12'd1900: rgb_data = 0;
12'd1901: rgb_data = 0;
12'd1902: rgb_data = 0;
12'd1903: rgb_data = 0;
12'd1904: rgb_data = 228;
12'd1905: rgb_data = 228;
12'd1906: rgb_data = 228;
12'd1907: rgb_data = 228;
12'd1908: rgb_data = 0;
12'd1909: rgb_data = 0;
12'd1910: rgb_data = 0;
12'd1911: rgb_data = 0;
12'd1912: rgb_data = 0;
12'd1913: rgb_data = 0;
12'd1914: rgb_data = 0;
12'd1915: rgb_data = 0;
12'd1916: rgb_data = 228;
12'd1917: rgb_data = 228;
12'd1918: rgb_data = 228;
12'd1919: rgb_data = 228;
12'd1920: rgb_data = 228;
12'd1921: rgb_data = 228;
12'd1922: rgb_data = 228;
12'd1923: rgb_data = 228;
12'd1924: rgb_data = 0;
12'd1925: rgb_data = 0;
12'd1926: rgb_data = 0;
12'd1927: rgb_data = 0;
12'd1928: rgb_data = 0;
12'd1929: rgb_data = 0;
12'd1930: rgb_data = 0;
12'd1931: rgb_data = 0;
12'd1932: rgb_data = 228;
12'd1933: rgb_data = 228;
12'd1934: rgb_data = 228;
12'd1935: rgb_data = 228;
12'd1936: rgb_data = 0;
12'd1937: rgb_data = 0;
12'd1938: rgb_data = 0;
12'd1939: rgb_data = 0;
12'd1940: rgb_data = 0;
12'd1941: rgb_data = 0;
12'd1942: rgb_data = 0;
12'd1943: rgb_data = 0;
12'd1944: rgb_data = 255;
12'd1945: rgb_data = 255;
12'd1946: rgb_data = 255;
12'd1947: rgb_data = 255;
12'd1948: rgb_data = 248;
12'd1949: rgb_data = 248;
12'd1950: rgb_data = 248;
12'd1951: rgb_data = 248;
12'd1952: rgb_data = 248;
12'd1953: rgb_data = 248;
12'd1954: rgb_data = 248;
12'd1955: rgb_data = 248;
12'd1956: rgb_data = 255;
12'd1957: rgb_data = 255;
12'd1958: rgb_data = 255;
12'd1959: rgb_data = 255;
12'd1960: rgb_data = 0;
12'd1961: rgb_data = 0;
12'd1962: rgb_data = 0;
12'd1963: rgb_data = 0;
12'd1964: rgb_data = 0;
12'd1965: rgb_data = 0;
12'd1966: rgb_data = 0;
12'd1967: rgb_data = 0;
12'd1968: rgb_data = 228;
12'd1969: rgb_data = 228;
12'd1970: rgb_data = 228;
12'd1971: rgb_data = 228;
12'd1972: rgb_data = 0;
12'd1973: rgb_data = 0;
12'd1974: rgb_data = 0;
12'd1975: rgb_data = 0;
12'd1976: rgb_data = 0;
12'd1977: rgb_data = 0;
12'd1978: rgb_data = 0;
12'd1979: rgb_data = 0;
12'd1980: rgb_data = 228;
12'd1981: rgb_data = 228;
12'd1982: rgb_data = 228;
12'd1983: rgb_data = 228;
12'd1984: rgb_data = 228;
12'd1985: rgb_data = 228;
12'd1986: rgb_data = 228;
12'd1987: rgb_data = 228;
12'd1988: rgb_data = 0;
12'd1989: rgb_data = 0;
12'd1990: rgb_data = 0;
12'd1991: rgb_data = 0;
12'd1992: rgb_data = 0;
12'd1993: rgb_data = 0;
12'd1994: rgb_data = 0;
12'd1995: rgb_data = 0;
12'd1996: rgb_data = 228;
12'd1997: rgb_data = 228;
12'd1998: rgb_data = 228;
12'd1999: rgb_data = 228;
12'd2000: rgb_data = 0;
12'd2001: rgb_data = 0;
12'd2002: rgb_data = 0;
12'd2003: rgb_data = 0;
12'd2004: rgb_data = 0;
12'd2005: rgb_data = 0;
12'd2006: rgb_data = 0;
12'd2007: rgb_data = 0;
12'd2008: rgb_data = 255;
12'd2009: rgb_data = 255;
12'd2010: rgb_data = 255;
12'd2011: rgb_data = 255;
12'd2012: rgb_data = 248;
12'd2013: rgb_data = 248;
12'd2014: rgb_data = 248;
12'd2015: rgb_data = 248;
12'd2016: rgb_data = 248;
12'd2017: rgb_data = 248;
12'd2018: rgb_data = 248;
12'd2019: rgb_data = 248;
12'd2020: rgb_data = 255;
12'd2021: rgb_data = 255;
12'd2022: rgb_data = 255;
12'd2023: rgb_data = 255;
12'd2024: rgb_data = 0;
12'd2025: rgb_data = 0;
12'd2026: rgb_data = 0;
12'd2027: rgb_data = 0;
12'd2028: rgb_data = 0;
12'd2029: rgb_data = 0;
12'd2030: rgb_data = 0;
12'd2031: rgb_data = 0;
12'd2032: rgb_data = 228;
12'd2033: rgb_data = 228;
12'd2034: rgb_data = 228;
12'd2035: rgb_data = 228;
12'd2036: rgb_data = 0;
12'd2037: rgb_data = 0;
12'd2038: rgb_data = 0;
12'd2039: rgb_data = 0;
12'd2040: rgb_data = 0;
12'd2041: rgb_data = 0;
12'd2042: rgb_data = 0;
12'd2043: rgb_data = 0;
12'd2044: rgb_data = 228;
12'd2045: rgb_data = 228;
12'd2046: rgb_data = 228;
12'd2047: rgb_data = 228;
12'd2048: rgb_data = 228;
12'd2049: rgb_data = 228;
12'd2050: rgb_data = 228;
12'd2051: rgb_data = 228;
12'd2052: rgb_data = 0;
12'd2053: rgb_data = 0;
12'd2054: rgb_data = 0;
12'd2055: rgb_data = 0;
12'd2056: rgb_data = 0;
12'd2057: rgb_data = 0;
12'd2058: rgb_data = 0;
12'd2059: rgb_data = 0;
12'd2060: rgb_data = 255;
12'd2061: rgb_data = 255;
12'd2062: rgb_data = 255;
12'd2063: rgb_data = 255;
12'd2064: rgb_data = 0;
12'd2065: rgb_data = 0;
12'd2066: rgb_data = 0;
12'd2067: rgb_data = 0;
12'd2068: rgb_data = 1;
12'd2069: rgb_data = 1;
12'd2070: rgb_data = 1;
12'd2071: rgb_data = 1;
12'd2072: rgb_data = 255;
12'd2073: rgb_data = 255;
12'd2074: rgb_data = 255;
12'd2075: rgb_data = 255;
12'd2076: rgb_data = 248;
12'd2077: rgb_data = 248;
12'd2078: rgb_data = 248;
12'd2079: rgb_data = 248;
12'd2080: rgb_data = 248;
12'd2081: rgb_data = 248;
12'd2082: rgb_data = 248;
12'd2083: rgb_data = 248;
12'd2084: rgb_data = 255;
12'd2085: rgb_data = 255;
12'd2086: rgb_data = 255;
12'd2087: rgb_data = 255;
12'd2088: rgb_data = 1;
12'd2089: rgb_data = 1;
12'd2090: rgb_data = 1;
12'd2091: rgb_data = 1;
12'd2092: rgb_data = 0;
12'd2093: rgb_data = 0;
12'd2094: rgb_data = 0;
12'd2095: rgb_data = 0;
12'd2096: rgb_data = 255;
12'd2097: rgb_data = 255;
12'd2098: rgb_data = 255;
12'd2099: rgb_data = 255;
12'd2100: rgb_data = 0;
12'd2101: rgb_data = 0;
12'd2102: rgb_data = 0;
12'd2103: rgb_data = 0;
12'd2104: rgb_data = 0;
12'd2105: rgb_data = 0;
12'd2106: rgb_data = 0;
12'd2107: rgb_data = 0;
12'd2108: rgb_data = 228;
12'd2109: rgb_data = 228;
12'd2110: rgb_data = 228;
12'd2111: rgb_data = 228;
12'd2112: rgb_data = 228;
12'd2113: rgb_data = 228;
12'd2114: rgb_data = 228;
12'd2115: rgb_data = 228;
12'd2116: rgb_data = 0;
12'd2117: rgb_data = 0;
12'd2118: rgb_data = 0;
12'd2119: rgb_data = 0;
12'd2120: rgb_data = 0;
12'd2121: rgb_data = 0;
12'd2122: rgb_data = 0;
12'd2123: rgb_data = 0;
12'd2124: rgb_data = 255;
12'd2125: rgb_data = 255;
12'd2126: rgb_data = 255;
12'd2127: rgb_data = 255;
12'd2128: rgb_data = 0;
12'd2129: rgb_data = 0;
12'd2130: rgb_data = 0;
12'd2131: rgb_data = 0;
12'd2132: rgb_data = 1;
12'd2133: rgb_data = 1;
12'd2134: rgb_data = 1;
12'd2135: rgb_data = 1;
12'd2136: rgb_data = 255;
12'd2137: rgb_data = 255;
12'd2138: rgb_data = 255;
12'd2139: rgb_data = 255;
12'd2140: rgb_data = 248;
12'd2141: rgb_data = 248;
12'd2142: rgb_data = 248;
12'd2143: rgb_data = 248;
12'd2144: rgb_data = 248;
12'd2145: rgb_data = 248;
12'd2146: rgb_data = 248;
12'd2147: rgb_data = 248;
12'd2148: rgb_data = 255;
12'd2149: rgb_data = 255;
12'd2150: rgb_data = 255;
12'd2151: rgb_data = 255;
12'd2152: rgb_data = 1;
12'd2153: rgb_data = 1;
12'd2154: rgb_data = 1;
12'd2155: rgb_data = 1;
12'd2156: rgb_data = 0;
12'd2157: rgb_data = 0;
12'd2158: rgb_data = 0;
12'd2159: rgb_data = 0;
12'd2160: rgb_data = 255;
12'd2161: rgb_data = 255;
12'd2162: rgb_data = 255;
12'd2163: rgb_data = 255;
12'd2164: rgb_data = 0;
12'd2165: rgb_data = 0;
12'd2166: rgb_data = 0;
12'd2167: rgb_data = 0;
12'd2168: rgb_data = 0;
12'd2169: rgb_data = 0;
12'd2170: rgb_data = 0;
12'd2171: rgb_data = 0;
12'd2172: rgb_data = 228;
12'd2173: rgb_data = 228;
12'd2174: rgb_data = 228;
12'd2175: rgb_data = 228;
12'd2176: rgb_data = 228;
12'd2177: rgb_data = 228;
12'd2178: rgb_data = 228;
12'd2179: rgb_data = 228;
12'd2180: rgb_data = 0;
12'd2181: rgb_data = 0;
12'd2182: rgb_data = 0;
12'd2183: rgb_data = 0;
12'd2184: rgb_data = 0;
12'd2185: rgb_data = 0;
12'd2186: rgb_data = 0;
12'd2187: rgb_data = 0;
12'd2188: rgb_data = 255;
12'd2189: rgb_data = 255;
12'd2190: rgb_data = 255;
12'd2191: rgb_data = 255;
12'd2192: rgb_data = 0;
12'd2193: rgb_data = 0;
12'd2194: rgb_data = 0;
12'd2195: rgb_data = 0;
12'd2196: rgb_data = 1;
12'd2197: rgb_data = 1;
12'd2198: rgb_data = 1;
12'd2199: rgb_data = 1;
12'd2200: rgb_data = 255;
12'd2201: rgb_data = 255;
12'd2202: rgb_data = 255;
12'd2203: rgb_data = 255;
12'd2204: rgb_data = 248;
12'd2205: rgb_data = 248;
12'd2206: rgb_data = 248;
12'd2207: rgb_data = 248;
12'd2208: rgb_data = 248;
12'd2209: rgb_data = 248;
12'd2210: rgb_data = 248;
12'd2211: rgb_data = 248;
12'd2212: rgb_data = 255;
12'd2213: rgb_data = 255;
12'd2214: rgb_data = 255;
12'd2215: rgb_data = 255;
12'd2216: rgb_data = 1;
12'd2217: rgb_data = 1;
12'd2218: rgb_data = 1;
12'd2219: rgb_data = 1;
12'd2220: rgb_data = 0;
12'd2221: rgb_data = 0;
12'd2222: rgb_data = 0;
12'd2223: rgb_data = 0;
12'd2224: rgb_data = 255;
12'd2225: rgb_data = 255;
12'd2226: rgb_data = 255;
12'd2227: rgb_data = 255;
12'd2228: rgb_data = 0;
12'd2229: rgb_data = 0;
12'd2230: rgb_data = 0;
12'd2231: rgb_data = 0;
12'd2232: rgb_data = 0;
12'd2233: rgb_data = 0;
12'd2234: rgb_data = 0;
12'd2235: rgb_data = 0;
12'd2236: rgb_data = 228;
12'd2237: rgb_data = 228;
12'd2238: rgb_data = 228;
12'd2239: rgb_data = 228;
12'd2240: rgb_data = 228;
12'd2241: rgb_data = 228;
12'd2242: rgb_data = 228;
12'd2243: rgb_data = 228;
12'd2244: rgb_data = 0;
12'd2245: rgb_data = 0;
12'd2246: rgb_data = 0;
12'd2247: rgb_data = 0;
12'd2248: rgb_data = 0;
12'd2249: rgb_data = 0;
12'd2250: rgb_data = 0;
12'd2251: rgb_data = 0;
12'd2252: rgb_data = 255;
12'd2253: rgb_data = 255;
12'd2254: rgb_data = 255;
12'd2255: rgb_data = 255;
12'd2256: rgb_data = 0;
12'd2257: rgb_data = 0;
12'd2258: rgb_data = 0;
12'd2259: rgb_data = 0;
12'd2260: rgb_data = 1;
12'd2261: rgb_data = 1;
12'd2262: rgb_data = 1;
12'd2263: rgb_data = 1;
12'd2264: rgb_data = 255;
12'd2265: rgb_data = 255;
12'd2266: rgb_data = 255;
12'd2267: rgb_data = 255;
12'd2268: rgb_data = 248;
12'd2269: rgb_data = 248;
12'd2270: rgb_data = 248;
12'd2271: rgb_data = 248;
12'd2272: rgb_data = 248;
12'd2273: rgb_data = 248;
12'd2274: rgb_data = 248;
12'd2275: rgb_data = 248;
12'd2276: rgb_data = 255;
12'd2277: rgb_data = 255;
12'd2278: rgb_data = 255;
12'd2279: rgb_data = 255;
12'd2280: rgb_data = 1;
12'd2281: rgb_data = 1;
12'd2282: rgb_data = 1;
12'd2283: rgb_data = 1;
12'd2284: rgb_data = 0;
12'd2285: rgb_data = 0;
12'd2286: rgb_data = 0;
12'd2287: rgb_data = 0;
12'd2288: rgb_data = 255;
12'd2289: rgb_data = 255;
12'd2290: rgb_data = 255;
12'd2291: rgb_data = 255;
12'd2292: rgb_data = 0;
12'd2293: rgb_data = 0;
12'd2294: rgb_data = 0;
12'd2295: rgb_data = 0;
12'd2296: rgb_data = 0;
12'd2297: rgb_data = 0;
12'd2298: rgb_data = 0;
12'd2299: rgb_data = 0;
12'd2300: rgb_data = 228;
12'd2301: rgb_data = 228;
12'd2302: rgb_data = 228;
12'd2303: rgb_data = 228;
12'd2304: rgb_data = 255;
12'd2305: rgb_data = 255;
12'd2306: rgb_data = 255;
12'd2307: rgb_data = 255;
12'd2308: rgb_data = 0;
12'd2309: rgb_data = 0;
12'd2310: rgb_data = 0;
12'd2311: rgb_data = 0;
12'd2312: rgb_data = 0;
12'd2313: rgb_data = 0;
12'd2314: rgb_data = 0;
12'd2315: rgb_data = 0;
12'd2316: rgb_data = 255;
12'd2317: rgb_data = 255;
12'd2318: rgb_data = 255;
12'd2319: rgb_data = 255;
12'd2320: rgb_data = 1;
12'd2321: rgb_data = 1;
12'd2322: rgb_data = 1;
12'd2323: rgb_data = 1;
12'd2324: rgb_data = 255;
12'd2325: rgb_data = 255;
12'd2326: rgb_data = 255;
12'd2327: rgb_data = 255;
12'd2328: rgb_data = 255;
12'd2329: rgb_data = 255;
12'd2330: rgb_data = 255;
12'd2331: rgb_data = 255;
12'd2332: rgb_data = 248;
12'd2333: rgb_data = 248;
12'd2334: rgb_data = 248;
12'd2335: rgb_data = 248;
12'd2336: rgb_data = 248;
12'd2337: rgb_data = 248;
12'd2338: rgb_data = 248;
12'd2339: rgb_data = 248;
12'd2340: rgb_data = 255;
12'd2341: rgb_data = 255;
12'd2342: rgb_data = 255;
12'd2343: rgb_data = 255;
12'd2344: rgb_data = 255;
12'd2345: rgb_data = 255;
12'd2346: rgb_data = 255;
12'd2347: rgb_data = 255;
12'd2348: rgb_data = 1;
12'd2349: rgb_data = 1;
12'd2350: rgb_data = 1;
12'd2351: rgb_data = 1;
12'd2352: rgb_data = 255;
12'd2353: rgb_data = 255;
12'd2354: rgb_data = 255;
12'd2355: rgb_data = 255;
12'd2356: rgb_data = 0;
12'd2357: rgb_data = 0;
12'd2358: rgb_data = 0;
12'd2359: rgb_data = 0;
12'd2360: rgb_data = 0;
12'd2361: rgb_data = 0;
12'd2362: rgb_data = 0;
12'd2363: rgb_data = 0;
12'd2364: rgb_data = 255;
12'd2365: rgb_data = 255;
12'd2366: rgb_data = 255;
12'd2367: rgb_data = 255;
12'd2368: rgb_data = 255;
12'd2369: rgb_data = 255;
12'd2370: rgb_data = 255;
12'd2371: rgb_data = 255;
12'd2372: rgb_data = 0;
12'd2373: rgb_data = 0;
12'd2374: rgb_data = 0;
12'd2375: rgb_data = 0;
12'd2376: rgb_data = 0;
12'd2377: rgb_data = 0;
12'd2378: rgb_data = 0;
12'd2379: rgb_data = 0;
12'd2380: rgb_data = 255;
12'd2381: rgb_data = 255;
12'd2382: rgb_data = 255;
12'd2383: rgb_data = 255;
12'd2384: rgb_data = 1;
12'd2385: rgb_data = 1;
12'd2386: rgb_data = 1;
12'd2387: rgb_data = 1;
12'd2388: rgb_data = 255;
12'd2389: rgb_data = 255;
12'd2390: rgb_data = 255;
12'd2391: rgb_data = 255;
12'd2392: rgb_data = 255;
12'd2393: rgb_data = 255;
12'd2394: rgb_data = 255;
12'd2395: rgb_data = 255;
12'd2396: rgb_data = 248;
12'd2397: rgb_data = 248;
12'd2398: rgb_data = 248;
12'd2399: rgb_data = 248;
12'd2400: rgb_data = 248;
12'd2401: rgb_data = 248;
12'd2402: rgb_data = 248;
12'd2403: rgb_data = 248;
12'd2404: rgb_data = 255;
12'd2405: rgb_data = 255;
12'd2406: rgb_data = 255;
12'd2407: rgb_data = 255;
12'd2408: rgb_data = 255;
12'd2409: rgb_data = 255;
12'd2410: rgb_data = 255;
12'd2411: rgb_data = 255;
12'd2412: rgb_data = 1;
12'd2413: rgb_data = 1;
12'd2414: rgb_data = 1;
12'd2415: rgb_data = 1;
12'd2416: rgb_data = 255;
12'd2417: rgb_data = 255;
12'd2418: rgb_data = 255;
12'd2419: rgb_data = 255;
12'd2420: rgb_data = 0;
12'd2421: rgb_data = 0;
12'd2422: rgb_data = 0;
12'd2423: rgb_data = 0;
12'd2424: rgb_data = 0;
12'd2425: rgb_data = 0;
12'd2426: rgb_data = 0;
12'd2427: rgb_data = 0;
12'd2428: rgb_data = 255;
12'd2429: rgb_data = 255;
12'd2430: rgb_data = 255;
12'd2431: rgb_data = 255;
12'd2432: rgb_data = 255;
12'd2433: rgb_data = 255;
12'd2434: rgb_data = 255;
12'd2435: rgb_data = 255;
12'd2436: rgb_data = 0;
12'd2437: rgb_data = 0;
12'd2438: rgb_data = 0;
12'd2439: rgb_data = 0;
12'd2440: rgb_data = 0;
12'd2441: rgb_data = 0;
12'd2442: rgb_data = 0;
12'd2443: rgb_data = 0;
12'd2444: rgb_data = 255;
12'd2445: rgb_data = 255;
12'd2446: rgb_data = 255;
12'd2447: rgb_data = 255;
12'd2448: rgb_data = 1;
12'd2449: rgb_data = 1;
12'd2450: rgb_data = 1;
12'd2451: rgb_data = 1;
12'd2452: rgb_data = 255;
12'd2453: rgb_data = 255;
12'd2454: rgb_data = 255;
12'd2455: rgb_data = 255;
12'd2456: rgb_data = 255;
12'd2457: rgb_data = 255;
12'd2458: rgb_data = 255;
12'd2459: rgb_data = 255;
12'd2460: rgb_data = 248;
12'd2461: rgb_data = 248;
12'd2462: rgb_data = 248;
12'd2463: rgb_data = 248;
12'd2464: rgb_data = 248;
12'd2465: rgb_data = 248;
12'd2466: rgb_data = 248;
12'd2467: rgb_data = 248;
12'd2468: rgb_data = 255;
12'd2469: rgb_data = 255;
12'd2470: rgb_data = 255;
12'd2471: rgb_data = 255;
12'd2472: rgb_data = 255;
12'd2473: rgb_data = 255;
12'd2474: rgb_data = 255;
12'd2475: rgb_data = 255;
12'd2476: rgb_data = 1;
12'd2477: rgb_data = 1;
12'd2478: rgb_data = 1;
12'd2479: rgb_data = 1;
12'd2480: rgb_data = 255;
12'd2481: rgb_data = 255;
12'd2482: rgb_data = 255;
12'd2483: rgb_data = 255;
12'd2484: rgb_data = 0;
12'd2485: rgb_data = 0;
12'd2486: rgb_data = 0;
12'd2487: rgb_data = 0;
12'd2488: rgb_data = 0;
12'd2489: rgb_data = 0;
12'd2490: rgb_data = 0;
12'd2491: rgb_data = 0;
12'd2492: rgb_data = 255;
12'd2493: rgb_data = 255;
12'd2494: rgb_data = 255;
12'd2495: rgb_data = 255;
12'd2496: rgb_data = 255;
12'd2497: rgb_data = 255;
12'd2498: rgb_data = 255;
12'd2499: rgb_data = 255;
12'd2500: rgb_data = 0;
12'd2501: rgb_data = 0;
12'd2502: rgb_data = 0;
12'd2503: rgb_data = 0;
12'd2504: rgb_data = 0;
12'd2505: rgb_data = 0;
12'd2506: rgb_data = 0;
12'd2507: rgb_data = 0;
12'd2508: rgb_data = 255;
12'd2509: rgb_data = 255;
12'd2510: rgb_data = 255;
12'd2511: rgb_data = 255;
12'd2512: rgb_data = 1;
12'd2513: rgb_data = 1;
12'd2514: rgb_data = 1;
12'd2515: rgb_data = 1;
12'd2516: rgb_data = 255;
12'd2517: rgb_data = 255;
12'd2518: rgb_data = 255;
12'd2519: rgb_data = 255;
12'd2520: rgb_data = 255;
12'd2521: rgb_data = 255;
12'd2522: rgb_data = 255;
12'd2523: rgb_data = 255;
12'd2524: rgb_data = 248;
12'd2525: rgb_data = 248;
12'd2526: rgb_data = 248;
12'd2527: rgb_data = 248;
12'd2528: rgb_data = 248;
12'd2529: rgb_data = 248;
12'd2530: rgb_data = 248;
12'd2531: rgb_data = 248;
12'd2532: rgb_data = 255;
12'd2533: rgb_data = 255;
12'd2534: rgb_data = 255;
12'd2535: rgb_data = 255;
12'd2536: rgb_data = 255;
12'd2537: rgb_data = 255;
12'd2538: rgb_data = 255;
12'd2539: rgb_data = 255;
12'd2540: rgb_data = 1;
12'd2541: rgb_data = 1;
12'd2542: rgb_data = 1;
12'd2543: rgb_data = 1;
12'd2544: rgb_data = 255;
12'd2545: rgb_data = 255;
12'd2546: rgb_data = 255;
12'd2547: rgb_data = 255;
12'd2548: rgb_data = 0;
12'd2549: rgb_data = 0;
12'd2550: rgb_data = 0;
12'd2551: rgb_data = 0;
12'd2552: rgb_data = 0;
12'd2553: rgb_data = 0;
12'd2554: rgb_data = 0;
12'd2555: rgb_data = 0;
12'd2556: rgb_data = 255;
12'd2557: rgb_data = 255;
12'd2558: rgb_data = 255;
12'd2559: rgb_data = 255;
12'd2560: rgb_data = 255;
12'd2561: rgb_data = 255;
12'd2562: rgb_data = 255;
12'd2563: rgb_data = 255;
12'd2564: rgb_data = 0;
12'd2565: rgb_data = 0;
12'd2566: rgb_data = 0;
12'd2567: rgb_data = 0;
12'd2568: rgb_data = 0;
12'd2569: rgb_data = 0;
12'd2570: rgb_data = 0;
12'd2571: rgb_data = 0;
12'd2572: rgb_data = 255;
12'd2573: rgb_data = 255;
12'd2574: rgb_data = 255;
12'd2575: rgb_data = 255;
12'd2576: rgb_data = 255;
12'd2577: rgb_data = 255;
12'd2578: rgb_data = 255;
12'd2579: rgb_data = 255;
12'd2580: rgb_data = 255;
12'd2581: rgb_data = 255;
12'd2582: rgb_data = 255;
12'd2583: rgb_data = 255;
12'd2584: rgb_data = 255;
12'd2585: rgb_data = 255;
12'd2586: rgb_data = 255;
12'd2587: rgb_data = 255;
12'd2588: rgb_data = 255;
12'd2589: rgb_data = 255;
12'd2590: rgb_data = 255;
12'd2591: rgb_data = 255;
12'd2592: rgb_data = 255;
12'd2593: rgb_data = 255;
12'd2594: rgb_data = 255;
12'd2595: rgb_data = 255;
12'd2596: rgb_data = 255;
12'd2597: rgb_data = 255;
12'd2598: rgb_data = 255;
12'd2599: rgb_data = 255;
12'd2600: rgb_data = 255;
12'd2601: rgb_data = 255;
12'd2602: rgb_data = 255;
12'd2603: rgb_data = 255;
12'd2604: rgb_data = 255;
12'd2605: rgb_data = 255;
12'd2606: rgb_data = 255;
12'd2607: rgb_data = 255;
12'd2608: rgb_data = 255;
12'd2609: rgb_data = 255;
12'd2610: rgb_data = 255;
12'd2611: rgb_data = 255;
12'd2612: rgb_data = 0;
12'd2613: rgb_data = 0;
12'd2614: rgb_data = 0;
12'd2615: rgb_data = 0;
12'd2616: rgb_data = 0;
12'd2617: rgb_data = 0;
12'd2618: rgb_data = 0;
12'd2619: rgb_data = 0;
12'd2620: rgb_data = 255;
12'd2621: rgb_data = 255;
12'd2622: rgb_data = 255;
12'd2623: rgb_data = 255;
12'd2624: rgb_data = 255;
12'd2625: rgb_data = 255;
12'd2626: rgb_data = 255;
12'd2627: rgb_data = 255;
12'd2628: rgb_data = 0;
12'd2629: rgb_data = 0;
12'd2630: rgb_data = 0;
12'd2631: rgb_data = 0;
12'd2632: rgb_data = 0;
12'd2633: rgb_data = 0;
12'd2634: rgb_data = 0;
12'd2635: rgb_data = 0;
12'd2636: rgb_data = 255;
12'd2637: rgb_data = 255;
12'd2638: rgb_data = 255;
12'd2639: rgb_data = 255;
12'd2640: rgb_data = 255;
12'd2641: rgb_data = 255;
12'd2642: rgb_data = 255;
12'd2643: rgb_data = 255;
12'd2644: rgb_data = 255;
12'd2645: rgb_data = 255;
12'd2646: rgb_data = 255;
12'd2647: rgb_data = 255;
12'd2648: rgb_data = 255;
12'd2649: rgb_data = 255;
12'd2650: rgb_data = 255;
12'd2651: rgb_data = 255;
12'd2652: rgb_data = 255;
12'd2653: rgb_data = 255;
12'd2654: rgb_data = 255;
12'd2655: rgb_data = 255;
12'd2656: rgb_data = 255;
12'd2657: rgb_data = 255;
12'd2658: rgb_data = 255;
12'd2659: rgb_data = 255;
12'd2660: rgb_data = 255;
12'd2661: rgb_data = 255;
12'd2662: rgb_data = 255;
12'd2663: rgb_data = 255;
12'd2664: rgb_data = 255;
12'd2665: rgb_data = 255;
12'd2666: rgb_data = 255;
12'd2667: rgb_data = 255;
12'd2668: rgb_data = 255;
12'd2669: rgb_data = 255;
12'd2670: rgb_data = 255;
12'd2671: rgb_data = 255;
12'd2672: rgb_data = 255;
12'd2673: rgb_data = 255;
12'd2674: rgb_data = 255;
12'd2675: rgb_data = 255;
12'd2676: rgb_data = 0;
12'd2677: rgb_data = 0;
12'd2678: rgb_data = 0;
12'd2679: rgb_data = 0;
12'd2680: rgb_data = 0;
12'd2681: rgb_data = 0;
12'd2682: rgb_data = 0;
12'd2683: rgb_data = 0;
12'd2684: rgb_data = 255;
12'd2685: rgb_data = 255;
12'd2686: rgb_data = 255;
12'd2687: rgb_data = 255;
12'd2688: rgb_data = 255;
12'd2689: rgb_data = 255;
12'd2690: rgb_data = 255;
12'd2691: rgb_data = 255;
12'd2692: rgb_data = 0;
12'd2693: rgb_data = 0;
12'd2694: rgb_data = 0;
12'd2695: rgb_data = 0;
12'd2696: rgb_data = 0;
12'd2697: rgb_data = 0;
12'd2698: rgb_data = 0;
12'd2699: rgb_data = 0;
12'd2700: rgb_data = 255;
12'd2701: rgb_data = 255;
12'd2702: rgb_data = 255;
12'd2703: rgb_data = 255;
12'd2704: rgb_data = 255;
12'd2705: rgb_data = 255;
12'd2706: rgb_data = 255;
12'd2707: rgb_data = 255;
12'd2708: rgb_data = 255;
12'd2709: rgb_data = 255;
12'd2710: rgb_data = 255;
12'd2711: rgb_data = 255;
12'd2712: rgb_data = 255;
12'd2713: rgb_data = 255;
12'd2714: rgb_data = 255;
12'd2715: rgb_data = 255;
12'd2716: rgb_data = 255;
12'd2717: rgb_data = 255;
12'd2718: rgb_data = 255;
12'd2719: rgb_data = 255;
12'd2720: rgb_data = 255;
12'd2721: rgb_data = 255;
12'd2722: rgb_data = 255;
12'd2723: rgb_data = 255;
12'd2724: rgb_data = 255;
12'd2725: rgb_data = 255;
12'd2726: rgb_data = 255;
12'd2727: rgb_data = 255;
12'd2728: rgb_data = 255;
12'd2729: rgb_data = 255;
12'd2730: rgb_data = 255;
12'd2731: rgb_data = 255;
12'd2732: rgb_data = 255;
12'd2733: rgb_data = 255;
12'd2734: rgb_data = 255;
12'd2735: rgb_data = 255;
12'd2736: rgb_data = 255;
12'd2737: rgb_data = 255;
12'd2738: rgb_data = 255;
12'd2739: rgb_data = 255;
12'd2740: rgb_data = 0;
12'd2741: rgb_data = 0;
12'd2742: rgb_data = 0;
12'd2743: rgb_data = 0;
12'd2744: rgb_data = 0;
12'd2745: rgb_data = 0;
12'd2746: rgb_data = 0;
12'd2747: rgb_data = 0;
12'd2748: rgb_data = 255;
12'd2749: rgb_data = 255;
12'd2750: rgb_data = 255;
12'd2751: rgb_data = 255;
12'd2752: rgb_data = 255;
12'd2753: rgb_data = 255;
12'd2754: rgb_data = 255;
12'd2755: rgb_data = 255;
12'd2756: rgb_data = 0;
12'd2757: rgb_data = 0;
12'd2758: rgb_data = 0;
12'd2759: rgb_data = 0;
12'd2760: rgb_data = 0;
12'd2761: rgb_data = 0;
12'd2762: rgb_data = 0;
12'd2763: rgb_data = 0;
12'd2764: rgb_data = 255;
12'd2765: rgb_data = 255;
12'd2766: rgb_data = 255;
12'd2767: rgb_data = 255;
12'd2768: rgb_data = 255;
12'd2769: rgb_data = 255;
12'd2770: rgb_data = 255;
12'd2771: rgb_data = 255;
12'd2772: rgb_data = 255;
12'd2773: rgb_data = 255;
12'd2774: rgb_data = 255;
12'd2775: rgb_data = 255;
12'd2776: rgb_data = 255;
12'd2777: rgb_data = 255;
12'd2778: rgb_data = 255;
12'd2779: rgb_data = 255;
12'd2780: rgb_data = 255;
12'd2781: rgb_data = 255;
12'd2782: rgb_data = 255;
12'd2783: rgb_data = 255;
12'd2784: rgb_data = 255;
12'd2785: rgb_data = 255;
12'd2786: rgb_data = 255;
12'd2787: rgb_data = 255;
12'd2788: rgb_data = 255;
12'd2789: rgb_data = 255;
12'd2790: rgb_data = 255;
12'd2791: rgb_data = 255;
12'd2792: rgb_data = 255;
12'd2793: rgb_data = 255;
12'd2794: rgb_data = 255;
12'd2795: rgb_data = 255;
12'd2796: rgb_data = 255;
12'd2797: rgb_data = 255;
12'd2798: rgb_data = 255;
12'd2799: rgb_data = 255;
12'd2800: rgb_data = 255;
12'd2801: rgb_data = 255;
12'd2802: rgb_data = 255;
12'd2803: rgb_data = 255;
12'd2804: rgb_data = 0;
12'd2805: rgb_data = 0;
12'd2806: rgb_data = 0;
12'd2807: rgb_data = 0;
12'd2808: rgb_data = 0;
12'd2809: rgb_data = 0;
12'd2810: rgb_data = 0;
12'd2811: rgb_data = 0;
12'd2812: rgb_data = 255;
12'd2813: rgb_data = 255;
12'd2814: rgb_data = 255;
12'd2815: rgb_data = 255;
12'd2816: rgb_data = 255;
12'd2817: rgb_data = 255;
12'd2818: rgb_data = 255;
12'd2819: rgb_data = 255;
12'd2820: rgb_data = 0;
12'd2821: rgb_data = 0;
12'd2822: rgb_data = 0;
12'd2823: rgb_data = 0;
12'd2824: rgb_data = 255;
12'd2825: rgb_data = 255;
12'd2826: rgb_data = 255;
12'd2827: rgb_data = 255;
12'd2828: rgb_data = 255;
12'd2829: rgb_data = 255;
12'd2830: rgb_data = 255;
12'd2831: rgb_data = 255;
12'd2832: rgb_data = 255;
12'd2833: rgb_data = 255;
12'd2834: rgb_data = 255;
12'd2835: rgb_data = 255;
12'd2836: rgb_data = 255;
12'd2837: rgb_data = 255;
12'd2838: rgb_data = 255;
12'd2839: rgb_data = 255;
12'd2840: rgb_data = 255;
12'd2841: rgb_data = 255;
12'd2842: rgb_data = 255;
12'd2843: rgb_data = 255;
12'd2844: rgb_data = 255;
12'd2845: rgb_data = 255;
12'd2846: rgb_data = 255;
12'd2847: rgb_data = 255;
12'd2848: rgb_data = 255;
12'd2849: rgb_data = 255;
12'd2850: rgb_data = 255;
12'd2851: rgb_data = 255;
12'd2852: rgb_data = 255;
12'd2853: rgb_data = 255;
12'd2854: rgb_data = 255;
12'd2855: rgb_data = 255;
12'd2856: rgb_data = 255;
12'd2857: rgb_data = 255;
12'd2858: rgb_data = 255;
12'd2859: rgb_data = 255;
12'd2860: rgb_data = 255;
12'd2861: rgb_data = 255;
12'd2862: rgb_data = 255;
12'd2863: rgb_data = 255;
12'd2864: rgb_data = 255;
12'd2865: rgb_data = 255;
12'd2866: rgb_data = 255;
12'd2867: rgb_data = 255;
12'd2868: rgb_data = 255;
12'd2869: rgb_data = 255;
12'd2870: rgb_data = 255;
12'd2871: rgb_data = 255;
12'd2872: rgb_data = 0;
12'd2873: rgb_data = 0;
12'd2874: rgb_data = 0;
12'd2875: rgb_data = 0;
12'd2876: rgb_data = 255;
12'd2877: rgb_data = 255;
12'd2878: rgb_data = 255;
12'd2879: rgb_data = 255;
12'd2880: rgb_data = 255;
12'd2881: rgb_data = 255;
12'd2882: rgb_data = 255;
12'd2883: rgb_data = 255;
12'd2884: rgb_data = 0;
12'd2885: rgb_data = 0;
12'd2886: rgb_data = 0;
12'd2887: rgb_data = 0;
12'd2888: rgb_data = 255;
12'd2889: rgb_data = 255;
12'd2890: rgb_data = 255;
12'd2891: rgb_data = 255;
12'd2892: rgb_data = 255;
12'd2893: rgb_data = 255;
12'd2894: rgb_data = 255;
12'd2895: rgb_data = 255;
12'd2896: rgb_data = 255;
12'd2897: rgb_data = 255;
12'd2898: rgb_data = 255;
12'd2899: rgb_data = 255;
12'd2900: rgb_data = 255;
12'd2901: rgb_data = 255;
12'd2902: rgb_data = 255;
12'd2903: rgb_data = 255;
12'd2904: rgb_data = 255;
12'd2905: rgb_data = 255;
12'd2906: rgb_data = 255;
12'd2907: rgb_data = 255;
12'd2908: rgb_data = 255;
12'd2909: rgb_data = 255;
12'd2910: rgb_data = 255;
12'd2911: rgb_data = 255;
12'd2912: rgb_data = 255;
12'd2913: rgb_data = 255;
12'd2914: rgb_data = 255;
12'd2915: rgb_data = 255;
12'd2916: rgb_data = 255;
12'd2917: rgb_data = 255;
12'd2918: rgb_data = 255;
12'd2919: rgb_data = 255;
12'd2920: rgb_data = 255;
12'd2921: rgb_data = 255;
12'd2922: rgb_data = 255;
12'd2923: rgb_data = 255;
12'd2924: rgb_data = 255;
12'd2925: rgb_data = 255;
12'd2926: rgb_data = 255;
12'd2927: rgb_data = 255;
12'd2928: rgb_data = 255;
12'd2929: rgb_data = 255;
12'd2930: rgb_data = 255;
12'd2931: rgb_data = 255;
12'd2932: rgb_data = 255;
12'd2933: rgb_data = 255;
12'd2934: rgb_data = 255;
12'd2935: rgb_data = 255;
12'd2936: rgb_data = 0;
12'd2937: rgb_data = 0;
12'd2938: rgb_data = 0;
12'd2939: rgb_data = 0;
12'd2940: rgb_data = 255;
12'd2941: rgb_data = 255;
12'd2942: rgb_data = 255;
12'd2943: rgb_data = 255;
12'd2944: rgb_data = 255;
12'd2945: rgb_data = 255;
12'd2946: rgb_data = 255;
12'd2947: rgb_data = 255;
12'd2948: rgb_data = 0;
12'd2949: rgb_data = 0;
12'd2950: rgb_data = 0;
12'd2951: rgb_data = 0;
12'd2952: rgb_data = 255;
12'd2953: rgb_data = 255;
12'd2954: rgb_data = 255;
12'd2955: rgb_data = 255;
12'd2956: rgb_data = 255;
12'd2957: rgb_data = 255;
12'd2958: rgb_data = 255;
12'd2959: rgb_data = 255;
12'd2960: rgb_data = 255;
12'd2961: rgb_data = 255;
12'd2962: rgb_data = 255;
12'd2963: rgb_data = 255;
12'd2964: rgb_data = 255;
12'd2965: rgb_data = 255;
12'd2966: rgb_data = 255;
12'd2967: rgb_data = 255;
12'd2968: rgb_data = 255;
12'd2969: rgb_data = 255;
12'd2970: rgb_data = 255;
12'd2971: rgb_data = 255;
12'd2972: rgb_data = 255;
12'd2973: rgb_data = 255;
12'd2974: rgb_data = 255;
12'd2975: rgb_data = 255;
12'd2976: rgb_data = 255;
12'd2977: rgb_data = 255;
12'd2978: rgb_data = 255;
12'd2979: rgb_data = 255;
12'd2980: rgb_data = 255;
12'd2981: rgb_data = 255;
12'd2982: rgb_data = 255;
12'd2983: rgb_data = 255;
12'd2984: rgb_data = 255;
12'd2985: rgb_data = 255;
12'd2986: rgb_data = 255;
12'd2987: rgb_data = 255;
12'd2988: rgb_data = 255;
12'd2989: rgb_data = 255;
12'd2990: rgb_data = 255;
12'd2991: rgb_data = 255;
12'd2992: rgb_data = 255;
12'd2993: rgb_data = 255;
12'd2994: rgb_data = 255;
12'd2995: rgb_data = 255;
12'd2996: rgb_data = 255;
12'd2997: rgb_data = 255;
12'd2998: rgb_data = 255;
12'd2999: rgb_data = 255;
12'd3000: rgb_data = 0;
12'd3001: rgb_data = 0;
12'd3002: rgb_data = 0;
12'd3003: rgb_data = 0;
12'd3004: rgb_data = 255;
12'd3005: rgb_data = 255;
12'd3006: rgb_data = 255;
12'd3007: rgb_data = 255;
12'd3008: rgb_data = 255;
12'd3009: rgb_data = 255;
12'd3010: rgb_data = 255;
12'd3011: rgb_data = 255;
12'd3012: rgb_data = 0;
12'd3013: rgb_data = 0;
12'd3014: rgb_data = 0;
12'd3015: rgb_data = 0;
12'd3016: rgb_data = 255;
12'd3017: rgb_data = 255;
12'd3018: rgb_data = 255;
12'd3019: rgb_data = 255;
12'd3020: rgb_data = 255;
12'd3021: rgb_data = 255;
12'd3022: rgb_data = 255;
12'd3023: rgb_data = 255;
12'd3024: rgb_data = 255;
12'd3025: rgb_data = 255;
12'd3026: rgb_data = 255;
12'd3027: rgb_data = 255;
12'd3028: rgb_data = 255;
12'd3029: rgb_data = 255;
12'd3030: rgb_data = 255;
12'd3031: rgb_data = 255;
12'd3032: rgb_data = 255;
12'd3033: rgb_data = 255;
12'd3034: rgb_data = 255;
12'd3035: rgb_data = 255;
12'd3036: rgb_data = 255;
12'd3037: rgb_data = 255;
12'd3038: rgb_data = 255;
12'd3039: rgb_data = 255;
12'd3040: rgb_data = 255;
12'd3041: rgb_data = 255;
12'd3042: rgb_data = 255;
12'd3043: rgb_data = 255;
12'd3044: rgb_data = 255;
12'd3045: rgb_data = 255;
12'd3046: rgb_data = 255;
12'd3047: rgb_data = 255;
12'd3048: rgb_data = 255;
12'd3049: rgb_data = 255;
12'd3050: rgb_data = 255;
12'd3051: rgb_data = 255;
12'd3052: rgb_data = 255;
12'd3053: rgb_data = 255;
12'd3054: rgb_data = 255;
12'd3055: rgb_data = 255;
12'd3056: rgb_data = 255;
12'd3057: rgb_data = 255;
12'd3058: rgb_data = 255;
12'd3059: rgb_data = 255;
12'd3060: rgb_data = 255;
12'd3061: rgb_data = 255;
12'd3062: rgb_data = 255;
12'd3063: rgb_data = 255;
12'd3064: rgb_data = 0;
12'd3065: rgb_data = 0;
12'd3066: rgb_data = 0;
12'd3067: rgb_data = 0;
12'd3068: rgb_data = 255;
12'd3069: rgb_data = 255;
12'd3070: rgb_data = 255;
12'd3071: rgb_data = 255;
12'd3072: rgb_data = 255;
12'd3073: rgb_data = 255;
12'd3074: rgb_data = 255;
12'd3075: rgb_data = 255;
12'd3076: rgb_data = 255;
12'd3077: rgb_data = 255;
12'd3078: rgb_data = 255;
12'd3079: rgb_data = 255;
12'd3080: rgb_data = 255;
12'd3081: rgb_data = 255;
12'd3082: rgb_data = 255;
12'd3083: rgb_data = 255;
12'd3084: rgb_data = 0;
12'd3085: rgb_data = 0;
12'd3086: rgb_data = 0;
12'd3087: rgb_data = 0;
12'd3088: rgb_data = 228;
12'd3089: rgb_data = 228;
12'd3090: rgb_data = 228;
12'd3091: rgb_data = 228;
12'd3092: rgb_data = 228;
12'd3093: rgb_data = 228;
12'd3094: rgb_data = 228;
12'd3095: rgb_data = 228;
12'd3096: rgb_data = 0;
12'd3097: rgb_data = 0;
12'd3098: rgb_data = 0;
12'd3099: rgb_data = 0;
12'd3100: rgb_data = 255;
12'd3101: rgb_data = 255;
12'd3102: rgb_data = 255;
12'd3103: rgb_data = 255;
12'd3104: rgb_data = 255;
12'd3105: rgb_data = 255;
12'd3106: rgb_data = 255;
12'd3107: rgb_data = 255;
12'd3108: rgb_data = 0;
12'd3109: rgb_data = 0;
12'd3110: rgb_data = 0;
12'd3111: rgb_data = 0;
12'd3112: rgb_data = 228;
12'd3113: rgb_data = 228;
12'd3114: rgb_data = 228;
12'd3115: rgb_data = 228;
12'd3116: rgb_data = 228;
12'd3117: rgb_data = 228;
12'd3118: rgb_data = 228;
12'd3119: rgb_data = 228;
12'd3120: rgb_data = 0;
12'd3121: rgb_data = 0;
12'd3122: rgb_data = 0;
12'd3123: rgb_data = 0;
12'd3124: rgb_data = 255;
12'd3125: rgb_data = 255;
12'd3126: rgb_data = 255;
12'd3127: rgb_data = 255;
12'd3128: rgb_data = 255;
12'd3129: rgb_data = 255;
12'd3130: rgb_data = 255;
12'd3131: rgb_data = 255;
12'd3132: rgb_data = 255;
12'd3133: rgb_data = 255;
12'd3134: rgb_data = 255;
12'd3135: rgb_data = 255;
12'd3136: rgb_data = 255;
12'd3137: rgb_data = 255;
12'd3138: rgb_data = 255;
12'd3139: rgb_data = 255;
12'd3140: rgb_data = 255;
12'd3141: rgb_data = 255;
12'd3142: rgb_data = 255;
12'd3143: rgb_data = 255;
12'd3144: rgb_data = 255;
12'd3145: rgb_data = 255;
12'd3146: rgb_data = 255;
12'd3147: rgb_data = 255;
12'd3148: rgb_data = 0;
12'd3149: rgb_data = 0;
12'd3150: rgb_data = 0;
12'd3151: rgb_data = 0;
12'd3152: rgb_data = 228;
12'd3153: rgb_data = 228;
12'd3154: rgb_data = 228;
12'd3155: rgb_data = 228;
12'd3156: rgb_data = 228;
12'd3157: rgb_data = 228;
12'd3158: rgb_data = 228;
12'd3159: rgb_data = 228;
12'd3160: rgb_data = 0;
12'd3161: rgb_data = 0;
12'd3162: rgb_data = 0;
12'd3163: rgb_data = 0;
12'd3164: rgb_data = 255;
12'd3165: rgb_data = 255;
12'd3166: rgb_data = 255;
12'd3167: rgb_data = 255;
12'd3168: rgb_data = 255;
12'd3169: rgb_data = 255;
12'd3170: rgb_data = 255;
12'd3171: rgb_data = 255;
12'd3172: rgb_data = 0;
12'd3173: rgb_data = 0;
12'd3174: rgb_data = 0;
12'd3175: rgb_data = 0;
12'd3176: rgb_data = 228;
12'd3177: rgb_data = 228;
12'd3178: rgb_data = 228;
12'd3179: rgb_data = 228;
12'd3180: rgb_data = 228;
12'd3181: rgb_data = 228;
12'd3182: rgb_data = 228;
12'd3183: rgb_data = 228;
12'd3184: rgb_data = 0;
12'd3185: rgb_data = 0;
12'd3186: rgb_data = 0;
12'd3187: rgb_data = 0;
12'd3188: rgb_data = 255;
12'd3189: rgb_data = 255;
12'd3190: rgb_data = 255;
12'd3191: rgb_data = 255;
12'd3192: rgb_data = 255;
12'd3193: rgb_data = 255;
12'd3194: rgb_data = 255;
12'd3195: rgb_data = 255;
12'd3196: rgb_data = 255;
12'd3197: rgb_data = 255;
12'd3198: rgb_data = 255;
12'd3199: rgb_data = 255;
12'd3200: rgb_data = 255;
12'd3201: rgb_data = 255;
12'd3202: rgb_data = 255;
12'd3203: rgb_data = 255;
12'd3204: rgb_data = 255;
12'd3205: rgb_data = 255;
12'd3206: rgb_data = 255;
12'd3207: rgb_data = 255;
12'd3208: rgb_data = 255;
12'd3209: rgb_data = 255;
12'd3210: rgb_data = 255;
12'd3211: rgb_data = 255;
12'd3212: rgb_data = 0;
12'd3213: rgb_data = 0;
12'd3214: rgb_data = 0;
12'd3215: rgb_data = 0;
12'd3216: rgb_data = 228;
12'd3217: rgb_data = 228;
12'd3218: rgb_data = 228;
12'd3219: rgb_data = 228;
12'd3220: rgb_data = 228;
12'd3221: rgb_data = 228;
12'd3222: rgb_data = 228;
12'd3223: rgb_data = 228;
12'd3224: rgb_data = 0;
12'd3225: rgb_data = 0;
12'd3226: rgb_data = 0;
12'd3227: rgb_data = 0;
12'd3228: rgb_data = 255;
12'd3229: rgb_data = 255;
12'd3230: rgb_data = 255;
12'd3231: rgb_data = 255;
12'd3232: rgb_data = 255;
12'd3233: rgb_data = 255;
12'd3234: rgb_data = 255;
12'd3235: rgb_data = 255;
12'd3236: rgb_data = 0;
12'd3237: rgb_data = 0;
12'd3238: rgb_data = 0;
12'd3239: rgb_data = 0;
12'd3240: rgb_data = 228;
12'd3241: rgb_data = 228;
12'd3242: rgb_data = 228;
12'd3243: rgb_data = 228;
12'd3244: rgb_data = 228;
12'd3245: rgb_data = 228;
12'd3246: rgb_data = 228;
12'd3247: rgb_data = 228;
12'd3248: rgb_data = 0;
12'd3249: rgb_data = 0;
12'd3250: rgb_data = 0;
12'd3251: rgb_data = 0;
12'd3252: rgb_data = 255;
12'd3253: rgb_data = 255;
12'd3254: rgb_data = 255;
12'd3255: rgb_data = 255;
12'd3256: rgb_data = 255;
12'd3257: rgb_data = 255;
12'd3258: rgb_data = 255;
12'd3259: rgb_data = 255;
12'd3260: rgb_data = 255;
12'd3261: rgb_data = 255;
12'd3262: rgb_data = 255;
12'd3263: rgb_data = 255;
12'd3264: rgb_data = 255;
12'd3265: rgb_data = 255;
12'd3266: rgb_data = 255;
12'd3267: rgb_data = 255;
12'd3268: rgb_data = 255;
12'd3269: rgb_data = 255;
12'd3270: rgb_data = 255;
12'd3271: rgb_data = 255;
12'd3272: rgb_data = 255;
12'd3273: rgb_data = 255;
12'd3274: rgb_data = 255;
12'd3275: rgb_data = 255;
12'd3276: rgb_data = 0;
12'd3277: rgb_data = 0;
12'd3278: rgb_data = 0;
12'd3279: rgb_data = 0;
12'd3280: rgb_data = 228;
12'd3281: rgb_data = 228;
12'd3282: rgb_data = 228;
12'd3283: rgb_data = 228;
12'd3284: rgb_data = 228;
12'd3285: rgb_data = 228;
12'd3286: rgb_data = 228;
12'd3287: rgb_data = 228;
12'd3288: rgb_data = 0;
12'd3289: rgb_data = 0;
12'd3290: rgb_data = 0;
12'd3291: rgb_data = 0;
12'd3292: rgb_data = 255;
12'd3293: rgb_data = 255;
12'd3294: rgb_data = 255;
12'd3295: rgb_data = 255;
12'd3296: rgb_data = 255;
12'd3297: rgb_data = 255;
12'd3298: rgb_data = 255;
12'd3299: rgb_data = 255;
12'd3300: rgb_data = 0;
12'd3301: rgb_data = 0;
12'd3302: rgb_data = 0;
12'd3303: rgb_data = 0;
12'd3304: rgb_data = 228;
12'd3305: rgb_data = 228;
12'd3306: rgb_data = 228;
12'd3307: rgb_data = 228;
12'd3308: rgb_data = 228;
12'd3309: rgb_data = 228;
12'd3310: rgb_data = 228;
12'd3311: rgb_data = 228;
12'd3312: rgb_data = 0;
12'd3313: rgb_data = 0;
12'd3314: rgb_data = 0;
12'd3315: rgb_data = 0;
12'd3316: rgb_data = 255;
12'd3317: rgb_data = 255;
12'd3318: rgb_data = 255;
12'd3319: rgb_data = 255;
12'd3320: rgb_data = 255;
12'd3321: rgb_data = 255;
12'd3322: rgb_data = 255;
12'd3323: rgb_data = 255;
12'd3324: rgb_data = 255;
12'd3325: rgb_data = 255;
12'd3326: rgb_data = 255;
12'd3327: rgb_data = 255;
12'd3328: rgb_data = 255;
12'd3329: rgb_data = 255;
12'd3330: rgb_data = 255;
12'd3331: rgb_data = 255;
12'd3332: rgb_data = 255;
12'd3333: rgb_data = 255;
12'd3334: rgb_data = 255;
12'd3335: rgb_data = 255;
12'd3336: rgb_data = 0;
12'd3337: rgb_data = 0;
12'd3338: rgb_data = 0;
12'd3339: rgb_data = 0;
12'd3340: rgb_data = 0;
12'd3341: rgb_data = 0;
12'd3342: rgb_data = 0;
12'd3343: rgb_data = 0;
12'd3344: rgb_data = 0;
12'd3345: rgb_data = 0;
12'd3346: rgb_data = 0;
12'd3347: rgb_data = 0;
12'd3348: rgb_data = 0;
12'd3349: rgb_data = 0;
12'd3350: rgb_data = 0;
12'd3351: rgb_data = 0;
12'd3352: rgb_data = 0;
12'd3353: rgb_data = 0;
12'd3354: rgb_data = 0;
12'd3355: rgb_data = 0;
12'd3356: rgb_data = 255;
12'd3357: rgb_data = 255;
12'd3358: rgb_data = 255;
12'd3359: rgb_data = 255;
12'd3360: rgb_data = 255;
12'd3361: rgb_data = 255;
12'd3362: rgb_data = 255;
12'd3363: rgb_data = 255;
12'd3364: rgb_data = 0;
12'd3365: rgb_data = 0;
12'd3366: rgb_data = 0;
12'd3367: rgb_data = 0;
12'd3368: rgb_data = 0;
12'd3369: rgb_data = 0;
12'd3370: rgb_data = 0;
12'd3371: rgb_data = 0;
12'd3372: rgb_data = 0;
12'd3373: rgb_data = 0;
12'd3374: rgb_data = 0;
12'd3375: rgb_data = 0;
12'd3376: rgb_data = 0;
12'd3377: rgb_data = 0;
12'd3378: rgb_data = 0;
12'd3379: rgb_data = 0;
12'd3380: rgb_data = 0;
12'd3381: rgb_data = 0;
12'd3382: rgb_data = 0;
12'd3383: rgb_data = 0;
12'd3384: rgb_data = 255;
12'd3385: rgb_data = 255;
12'd3386: rgb_data = 255;
12'd3387: rgb_data = 255;
12'd3388: rgb_data = 255;
12'd3389: rgb_data = 255;
12'd3390: rgb_data = 255;
12'd3391: rgb_data = 255;
12'd3392: rgb_data = 255;
12'd3393: rgb_data = 255;
12'd3394: rgb_data = 255;
12'd3395: rgb_data = 255;
12'd3396: rgb_data = 255;
12'd3397: rgb_data = 255;
12'd3398: rgb_data = 255;
12'd3399: rgb_data = 255;
12'd3400: rgb_data = 0;
12'd3401: rgb_data = 0;
12'd3402: rgb_data = 0;
12'd3403: rgb_data = 0;
12'd3404: rgb_data = 0;
12'd3405: rgb_data = 0;
12'd3406: rgb_data = 0;
12'd3407: rgb_data = 0;
12'd3408: rgb_data = 0;
12'd3409: rgb_data = 0;
12'd3410: rgb_data = 0;
12'd3411: rgb_data = 0;
12'd3412: rgb_data = 0;
12'd3413: rgb_data = 0;
12'd3414: rgb_data = 0;
12'd3415: rgb_data = 0;
12'd3416: rgb_data = 0;
12'd3417: rgb_data = 0;
12'd3418: rgb_data = 0;
12'd3419: rgb_data = 0;
12'd3420: rgb_data = 255;
12'd3421: rgb_data = 255;
12'd3422: rgb_data = 255;
12'd3423: rgb_data = 255;
12'd3424: rgb_data = 255;
12'd3425: rgb_data = 255;
12'd3426: rgb_data = 255;
12'd3427: rgb_data = 255;
12'd3428: rgb_data = 0;
12'd3429: rgb_data = 0;
12'd3430: rgb_data = 0;
12'd3431: rgb_data = 0;
12'd3432: rgb_data = 0;
12'd3433: rgb_data = 0;
12'd3434: rgb_data = 0;
12'd3435: rgb_data = 0;
12'd3436: rgb_data = 0;
12'd3437: rgb_data = 0;
12'd3438: rgb_data = 0;
12'd3439: rgb_data = 0;
12'd3440: rgb_data = 0;
12'd3441: rgb_data = 0;
12'd3442: rgb_data = 0;
12'd3443: rgb_data = 0;
12'd3444: rgb_data = 0;
12'd3445: rgb_data = 0;
12'd3446: rgb_data = 0;
12'd3447: rgb_data = 0;
12'd3448: rgb_data = 255;
12'd3449: rgb_data = 255;
12'd3450: rgb_data = 255;
12'd3451: rgb_data = 255;
12'd3452: rgb_data = 255;
12'd3453: rgb_data = 255;
12'd3454: rgb_data = 255;
12'd3455: rgb_data = 255;
12'd3456: rgb_data = 255;
12'd3457: rgb_data = 255;
12'd3458: rgb_data = 255;
12'd3459: rgb_data = 255;
12'd3460: rgb_data = 255;
12'd3461: rgb_data = 255;
12'd3462: rgb_data = 255;
12'd3463: rgb_data = 255;
12'd3464: rgb_data = 0;
12'd3465: rgb_data = 0;
12'd3466: rgb_data = 0;
12'd3467: rgb_data = 0;
12'd3468: rgb_data = 0;
12'd3469: rgb_data = 0;
12'd3470: rgb_data = 0;
12'd3471: rgb_data = 0;
12'd3472: rgb_data = 0;
12'd3473: rgb_data = 0;
12'd3474: rgb_data = 0;
12'd3475: rgb_data = 0;
12'd3476: rgb_data = 0;
12'd3477: rgb_data = 0;
12'd3478: rgb_data = 0;
12'd3479: rgb_data = 0;
12'd3480: rgb_data = 0;
12'd3481: rgb_data = 0;
12'd3482: rgb_data = 0;
12'd3483: rgb_data = 0;
12'd3484: rgb_data = 255;
12'd3485: rgb_data = 255;
12'd3486: rgb_data = 255;
12'd3487: rgb_data = 255;
12'd3488: rgb_data = 255;
12'd3489: rgb_data = 255;
12'd3490: rgb_data = 255;
12'd3491: rgb_data = 255;
12'd3492: rgb_data = 0;
12'd3493: rgb_data = 0;
12'd3494: rgb_data = 0;
12'd3495: rgb_data = 0;
12'd3496: rgb_data = 0;
12'd3497: rgb_data = 0;
12'd3498: rgb_data = 0;
12'd3499: rgb_data = 0;
12'd3500: rgb_data = 0;
12'd3501: rgb_data = 0;
12'd3502: rgb_data = 0;
12'd3503: rgb_data = 0;
12'd3504: rgb_data = 0;
12'd3505: rgb_data = 0;
12'd3506: rgb_data = 0;
12'd3507: rgb_data = 0;
12'd3508: rgb_data = 0;
12'd3509: rgb_data = 0;
12'd3510: rgb_data = 0;
12'd3511: rgb_data = 0;
12'd3512: rgb_data = 255;
12'd3513: rgb_data = 255;
12'd3514: rgb_data = 255;
12'd3515: rgb_data = 255;
12'd3516: rgb_data = 255;
12'd3517: rgb_data = 255;
12'd3518: rgb_data = 255;
12'd3519: rgb_data = 255;
12'd3520: rgb_data = 255;
12'd3521: rgb_data = 255;
12'd3522: rgb_data = 255;
12'd3523: rgb_data = 255;
12'd3524: rgb_data = 255;
12'd3525: rgb_data = 255;
12'd3526: rgb_data = 255;
12'd3527: rgb_data = 255;
12'd3528: rgb_data = 0;
12'd3529: rgb_data = 0;
12'd3530: rgb_data = 0;
12'd3531: rgb_data = 0;
12'd3532: rgb_data = 0;
12'd3533: rgb_data = 0;
12'd3534: rgb_data = 0;
12'd3535: rgb_data = 0;
12'd3536: rgb_data = 0;
12'd3537: rgb_data = 0;
12'd3538: rgb_data = 0;
12'd3539: rgb_data = 0;
12'd3540: rgb_data = 0;
12'd3541: rgb_data = 0;
12'd3542: rgb_data = 0;
12'd3543: rgb_data = 0;
12'd3544: rgb_data = 0;
12'd3545: rgb_data = 0;
12'd3546: rgb_data = 0;
12'd3547: rgb_data = 0;
12'd3548: rgb_data = 255;
12'd3549: rgb_data = 255;
12'd3550: rgb_data = 255;
12'd3551: rgb_data = 255;
12'd3552: rgb_data = 255;
12'd3553: rgb_data = 255;
12'd3554: rgb_data = 255;
12'd3555: rgb_data = 255;
12'd3556: rgb_data = 0;
12'd3557: rgb_data = 0;
12'd3558: rgb_data = 0;
12'd3559: rgb_data = 0;
12'd3560: rgb_data = 0;
12'd3561: rgb_data = 0;
12'd3562: rgb_data = 0;
12'd3563: rgb_data = 0;
12'd3564: rgb_data = 0;
12'd3565: rgb_data = 0;
12'd3566: rgb_data = 0;
12'd3567: rgb_data = 0;
12'd3568: rgb_data = 0;
12'd3569: rgb_data = 0;
12'd3570: rgb_data = 0;
12'd3571: rgb_data = 0;
12'd3572: rgb_data = 0;
12'd3573: rgb_data = 0;
12'd3574: rgb_data = 0;
12'd3575: rgb_data = 0;
12'd3576: rgb_data = 255;
12'd3577: rgb_data = 255;
12'd3578: rgb_data = 255;
12'd3579: rgb_data = 255;
12'd3580: rgb_data = 255;
12'd3581: rgb_data = 255;
12'd3582: rgb_data = 255;
12'd3583: rgb_data = 255;
12'd3584: rgb_data = 0;
12'd3585: rgb_data = 0;
12'd3586: rgb_data = 0;
12'd3587: rgb_data = 0;
12'd3588: rgb_data = 0;
12'd3589: rgb_data = 0;
12'd3590: rgb_data = 0;
12'd3591: rgb_data = 0;
12'd3592: rgb_data = 0;
12'd3593: rgb_data = 0;
12'd3594: rgb_data = 0;
12'd3595: rgb_data = 0;
12'd3596: rgb_data = 0;
12'd3597: rgb_data = 0;
12'd3598: rgb_data = 0;
12'd3599: rgb_data = 0;
12'd3600: rgb_data = 0;
12'd3601: rgb_data = 0;
12'd3602: rgb_data = 0;
12'd3603: rgb_data = 0;
12'd3604: rgb_data = 0;
12'd3605: rgb_data = 0;
12'd3606: rgb_data = 0;
12'd3607: rgb_data = 0;
12'd3608: rgb_data = 0;
12'd3609: rgb_data = 0;
12'd3610: rgb_data = 0;
12'd3611: rgb_data = 0;
12'd3612: rgb_data = 0;
12'd3613: rgb_data = 0;
12'd3614: rgb_data = 0;
12'd3615: rgb_data = 0;
12'd3616: rgb_data = 0;
12'd3617: rgb_data = 0;
12'd3618: rgb_data = 0;
12'd3619: rgb_data = 0;
12'd3620: rgb_data = 0;
12'd3621: rgb_data = 0;
12'd3622: rgb_data = 0;
12'd3623: rgb_data = 0;
12'd3624: rgb_data = 0;
12'd3625: rgb_data = 0;
12'd3626: rgb_data = 0;
12'd3627: rgb_data = 0;
12'd3628: rgb_data = 0;
12'd3629: rgb_data = 0;
12'd3630: rgb_data = 0;
12'd3631: rgb_data = 0;
12'd3632: rgb_data = 0;
12'd3633: rgb_data = 0;
12'd3634: rgb_data = 0;
12'd3635: rgb_data = 0;
12'd3636: rgb_data = 0;
12'd3637: rgb_data = 0;
12'd3638: rgb_data = 0;
12'd3639: rgb_data = 0;
12'd3640: rgb_data = 0;
12'd3641: rgb_data = 0;
12'd3642: rgb_data = 0;
12'd3643: rgb_data = 0;
12'd3644: rgb_data = 0;
12'd3645: rgb_data = 0;
12'd3646: rgb_data = 0;
12'd3647: rgb_data = 0;
12'd3648: rgb_data = 0;
12'd3649: rgb_data = 0;
12'd3650: rgb_data = 0;
12'd3651: rgb_data = 0;
12'd3652: rgb_data = 0;
12'd3653: rgb_data = 0;
12'd3654: rgb_data = 0;
12'd3655: rgb_data = 0;
12'd3656: rgb_data = 0;
12'd3657: rgb_data = 0;
12'd3658: rgb_data = 0;
12'd3659: rgb_data = 0;
12'd3660: rgb_data = 0;
12'd3661: rgb_data = 0;
12'd3662: rgb_data = 0;
12'd3663: rgb_data = 0;
12'd3664: rgb_data = 0;
12'd3665: rgb_data = 0;
12'd3666: rgb_data = 0;
12'd3667: rgb_data = 0;
12'd3668: rgb_data = 0;
12'd3669: rgb_data = 0;
12'd3670: rgb_data = 0;
12'd3671: rgb_data = 0;
12'd3672: rgb_data = 0;
12'd3673: rgb_data = 0;
12'd3674: rgb_data = 0;
12'd3675: rgb_data = 0;
12'd3676: rgb_data = 0;
12'd3677: rgb_data = 0;
12'd3678: rgb_data = 0;
12'd3679: rgb_data = 0;
12'd3680: rgb_data = 0;
12'd3681: rgb_data = 0;
12'd3682: rgb_data = 0;
12'd3683: rgb_data = 0;
12'd3684: rgb_data = 0;
12'd3685: rgb_data = 0;
12'd3686: rgb_data = 0;
12'd3687: rgb_data = 0;
12'd3688: rgb_data = 0;
12'd3689: rgb_data = 0;
12'd3690: rgb_data = 0;
12'd3691: rgb_data = 0;
12'd3692: rgb_data = 0;
12'd3693: rgb_data = 0;
12'd3694: rgb_data = 0;
12'd3695: rgb_data = 0;
12'd3696: rgb_data = 0;
12'd3697: rgb_data = 0;
12'd3698: rgb_data = 0;
12'd3699: rgb_data = 0;
12'd3700: rgb_data = 0;
12'd3701: rgb_data = 0;
12'd3702: rgb_data = 0;
12'd3703: rgb_data = 0;
12'd3704: rgb_data = 0;
12'd3705: rgb_data = 0;
12'd3706: rgb_data = 0;
12'd3707: rgb_data = 0;
12'd3708: rgb_data = 0;
12'd3709: rgb_data = 0;
12'd3710: rgb_data = 0;
12'd3711: rgb_data = 0;
12'd3712: rgb_data = 0;
12'd3713: rgb_data = 0;
12'd3714: rgb_data = 0;
12'd3715: rgb_data = 0;
12'd3716: rgb_data = 0;
12'd3717: rgb_data = 0;
12'd3718: rgb_data = 0;
12'd3719: rgb_data = 0;
12'd3720: rgb_data = 0;
12'd3721: rgb_data = 0;
12'd3722: rgb_data = 0;
12'd3723: rgb_data = 0;
12'd3724: rgb_data = 0;
12'd3725: rgb_data = 0;
12'd3726: rgb_data = 0;
12'd3727: rgb_data = 0;
12'd3728: rgb_data = 0;
12'd3729: rgb_data = 0;
12'd3730: rgb_data = 0;
12'd3731: rgb_data = 0;
12'd3732: rgb_data = 0;
12'd3733: rgb_data = 0;
12'd3734: rgb_data = 0;
12'd3735: rgb_data = 0;
12'd3736: rgb_data = 0;
12'd3737: rgb_data = 0;
12'd3738: rgb_data = 0;
12'd3739: rgb_data = 0;
12'd3740: rgb_data = 0;
12'd3741: rgb_data = 0;
12'd3742: rgb_data = 0;
12'd3743: rgb_data = 0;
12'd3744: rgb_data = 0;
12'd3745: rgb_data = 0;
12'd3746: rgb_data = 0;
12'd3747: rgb_data = 0;
12'd3748: rgb_data = 0;
12'd3749: rgb_data = 0;
12'd3750: rgb_data = 0;
12'd3751: rgb_data = 0;
12'd3752: rgb_data = 0;
12'd3753: rgb_data = 0;
12'd3754: rgb_data = 0;
12'd3755: rgb_data = 0;
12'd3756: rgb_data = 0;
12'd3757: rgb_data = 0;
12'd3758: rgb_data = 0;
12'd3759: rgb_data = 0;
12'd3760: rgb_data = 0;
12'd3761: rgb_data = 0;
12'd3762: rgb_data = 0;
12'd3763: rgb_data = 0;
12'd3764: rgb_data = 0;
12'd3765: rgb_data = 0;
12'd3766: rgb_data = 0;
12'd3767: rgb_data = 0;
12'd3768: rgb_data = 0;
12'd3769: rgb_data = 0;
12'd3770: rgb_data = 0;
12'd3771: rgb_data = 0;
12'd3772: rgb_data = 0;
12'd3773: rgb_data = 0;
12'd3774: rgb_data = 0;
12'd3775: rgb_data = 0;
12'd3776: rgb_data = 0;
12'd3777: rgb_data = 0;
12'd3778: rgb_data = 0;
12'd3779: rgb_data = 0;
12'd3780: rgb_data = 0;
12'd3781: rgb_data = 0;
12'd3782: rgb_data = 0;
12'd3783: rgb_data = 0;
12'd3784: rgb_data = 0;
12'd3785: rgb_data = 0;
12'd3786: rgb_data = 0;
12'd3787: rgb_data = 0;
12'd3788: rgb_data = 0;
12'd3789: rgb_data = 0;
12'd3790: rgb_data = 0;
12'd3791: rgb_data = 0;
12'd3792: rgb_data = 0;
12'd3793: rgb_data = 0;
12'd3794: rgb_data = 0;
12'd3795: rgb_data = 0;
12'd3796: rgb_data = 0;
12'd3797: rgb_data = 0;
12'd3798: rgb_data = 0;
12'd3799: rgb_data = 0;
12'd3800: rgb_data = 0;
12'd3801: rgb_data = 0;
12'd3802: rgb_data = 0;
12'd3803: rgb_data = 0;
12'd3804: rgb_data = 0;
12'd3805: rgb_data = 0;
12'd3806: rgb_data = 0;
12'd3807: rgb_data = 0;
12'd3808: rgb_data = 0;
12'd3809: rgb_data = 0;
12'd3810: rgb_data = 0;
12'd3811: rgb_data = 0;
12'd3812: rgb_data = 0;
12'd3813: rgb_data = 0;
12'd3814: rgb_data = 0;
12'd3815: rgb_data = 0;
12'd3816: rgb_data = 0;
12'd3817: rgb_data = 0;
12'd3818: rgb_data = 0;
12'd3819: rgb_data = 0;
12'd3820: rgb_data = 0;
12'd3821: rgb_data = 0;
12'd3822: rgb_data = 0;
12'd3823: rgb_data = 0;
12'd3824: rgb_data = 0;
12'd3825: rgb_data = 0;
12'd3826: rgb_data = 0;
12'd3827: rgb_data = 0;
12'd3828: rgb_data = 0;
12'd3829: rgb_data = 0;
12'd3830: rgb_data = 0;
12'd3831: rgb_data = 0;
12'd3832: rgb_data = 0;
12'd3833: rgb_data = 0;
12'd3834: rgb_data = 0;
12'd3835: rgb_data = 0;
12'd3836: rgb_data = 0;
12'd3837: rgb_data = 0;
12'd3838: rgb_data = 0;
12'd3839: rgb_data = 0;
12'd3840: rgb_data = 0;
12'd3841: rgb_data = 0;
12'd3842: rgb_data = 0;
12'd3843: rgb_data = 0;
12'd3844: rgb_data = 0;
12'd3845: rgb_data = 0;
12'd3846: rgb_data = 0;
12'd3847: rgb_data = 0;
12'd3848: rgb_data = 0;
12'd3849: rgb_data = 0;
12'd3850: rgb_data = 0;
12'd3851: rgb_data = 0;
12'd3852: rgb_data = 0;
12'd3853: rgb_data = 0;
12'd3854: rgb_data = 0;
12'd3855: rgb_data = 0;
12'd3856: rgb_data = 0;
12'd3857: rgb_data = 0;
12'd3858: rgb_data = 0;
12'd3859: rgb_data = 0;
12'd3860: rgb_data = 0;
12'd3861: rgb_data = 0;
12'd3862: rgb_data = 0;
12'd3863: rgb_data = 0;
12'd3864: rgb_data = 0;
12'd3865: rgb_data = 0;
12'd3866: rgb_data = 0;
12'd3867: rgb_data = 0;
12'd3868: rgb_data = 0;
12'd3869: rgb_data = 0;
12'd3870: rgb_data = 0;
12'd3871: rgb_data = 0;
12'd3872: rgb_data = 0;
12'd3873: rgb_data = 0;
12'd3874: rgb_data = 0;
12'd3875: rgb_data = 0;
12'd3876: rgb_data = 0;
12'd3877: rgb_data = 0;
12'd3878: rgb_data = 0;
12'd3879: rgb_data = 0;
12'd3880: rgb_data = 0;
12'd3881: rgb_data = 0;
12'd3882: rgb_data = 0;
12'd3883: rgb_data = 0;
12'd3884: rgb_data = 0;
12'd3885: rgb_data = 0;
12'd3886: rgb_data = 0;
12'd3887: rgb_data = 0;
12'd3888: rgb_data = 0;
12'd3889: rgb_data = 0;
12'd3890: rgb_data = 0;
12'd3891: rgb_data = 0;
12'd3892: rgb_data = 0;
12'd3893: rgb_data = 0;
12'd3894: rgb_data = 0;
12'd3895: rgb_data = 0;
12'd3896: rgb_data = 0;
12'd3897: rgb_data = 0;
12'd3898: rgb_data = 0;
12'd3899: rgb_data = 0;
12'd3900: rgb_data = 0;
12'd3901: rgb_data = 0;
12'd3902: rgb_data = 0;
12'd3903: rgb_data = 0;
12'd3904: rgb_data = 0;
12'd3905: rgb_data = 0;
12'd3906: rgb_data = 0;
12'd3907: rgb_data = 0;
12'd3908: rgb_data = 0;
12'd3909: rgb_data = 0;
12'd3910: rgb_data = 0;
12'd3911: rgb_data = 0;
12'd3912: rgb_data = 0;
12'd3913: rgb_data = 0;
12'd3914: rgb_data = 0;
12'd3915: rgb_data = 0;
12'd3916: rgb_data = 0;
12'd3917: rgb_data = 0;
12'd3918: rgb_data = 0;
12'd3919: rgb_data = 0;
12'd3920: rgb_data = 0;
12'd3921: rgb_data = 0;
12'd3922: rgb_data = 0;
12'd3923: rgb_data = 0;
12'd3924: rgb_data = 0;
12'd3925: rgb_data = 0;
12'd3926: rgb_data = 0;
12'd3927: rgb_data = 0;
12'd3928: rgb_data = 0;
12'd3929: rgb_data = 0;
12'd3930: rgb_data = 0;
12'd3931: rgb_data = 0;
12'd3932: rgb_data = 0;
12'd3933: rgb_data = 0;
12'd3934: rgb_data = 0;
12'd3935: rgb_data = 0;
12'd3936: rgb_data = 0;
12'd3937: rgb_data = 0;
12'd3938: rgb_data = 0;
12'd3939: rgb_data = 0;
12'd3940: rgb_data = 0;
12'd3941: rgb_data = 0;
12'd3942: rgb_data = 0;
12'd3943: rgb_data = 0;
12'd3944: rgb_data = 0;
12'd3945: rgb_data = 0;
12'd3946: rgb_data = 0;
12'd3947: rgb_data = 0;
12'd3948: rgb_data = 0;
12'd3949: rgb_data = 0;
12'd3950: rgb_data = 0;
12'd3951: rgb_data = 0;
12'd3952: rgb_data = 0;
12'd3953: rgb_data = 0;
12'd3954: rgb_data = 0;
12'd3955: rgb_data = 0;
12'd3956: rgb_data = 0;
12'd3957: rgb_data = 0;
12'd3958: rgb_data = 0;
12'd3959: rgb_data = 0;
12'd3960: rgb_data = 0;
12'd3961: rgb_data = 0;
12'd3962: rgb_data = 0;
12'd3963: rgb_data = 0;
12'd3964: rgb_data = 0;
12'd3965: rgb_data = 0;
12'd3966: rgb_data = 0;
12'd3967: rgb_data = 0;
12'd3968: rgb_data = 0;
12'd3969: rgb_data = 0;
12'd3970: rgb_data = 0;
12'd3971: rgb_data = 0;
12'd3972: rgb_data = 0;
12'd3973: rgb_data = 0;
12'd3974: rgb_data = 0;
12'd3975: rgb_data = 0;
12'd3976: rgb_data = 0;
12'd3977: rgb_data = 0;
12'd3978: rgb_data = 0;
12'd3979: rgb_data = 0;
12'd3980: rgb_data = 0;
12'd3981: rgb_data = 0;
12'd3982: rgb_data = 0;
12'd3983: rgb_data = 0;
12'd3984: rgb_data = 0;
12'd3985: rgb_data = 0;
12'd3986: rgb_data = 0;
12'd3987: rgb_data = 0;
12'd3988: rgb_data = 0;
12'd3989: rgb_data = 0;
12'd3990: rgb_data = 0;
12'd3991: rgb_data = 0;
12'd3992: rgb_data = 0;
12'd3993: rgb_data = 0;
12'd3994: rgb_data = 0;
12'd3995: rgb_data = 0;
12'd3996: rgb_data = 0;
12'd3997: rgb_data = 0;
12'd3998: rgb_data = 0;
12'd3999: rgb_data = 0;
12'd4000: rgb_data = 0;
12'd4001: rgb_data = 0;
12'd4002: rgb_data = 0;
12'd4003: rgb_data = 0;
12'd4004: rgb_data = 0;
12'd4005: rgb_data = 0;
12'd4006: rgb_data = 0;
12'd4007: rgb_data = 0;
12'd4008: rgb_data = 0;
12'd4009: rgb_data = 0;
12'd4010: rgb_data = 0;
12'd4011: rgb_data = 0;
12'd4012: rgb_data = 0;
12'd4013: rgb_data = 0;
12'd4014: rgb_data = 0;
12'd4015: rgb_data = 0;
12'd4016: rgb_data = 0;
12'd4017: rgb_data = 0;
12'd4018: rgb_data = 0;
12'd4019: rgb_data = 0;
12'd4020: rgb_data = 0;
12'd4021: rgb_data = 0;
12'd4022: rgb_data = 0;
12'd4023: rgb_data = 0;
12'd4024: rgb_data = 0;
12'd4025: rgb_data = 0;
12'd4026: rgb_data = 0;
12'd4027: rgb_data = 0;
12'd4028: rgb_data = 0;
12'd4029: rgb_data = 0;
12'd4030: rgb_data = 0;
12'd4031: rgb_data = 0;
12'd4032: rgb_data = 0;
12'd4033: rgb_data = 0;
12'd4034: rgb_data = 0;
12'd4035: rgb_data = 0;
12'd4036: rgb_data = 0;
12'd4037: rgb_data = 0;
12'd4038: rgb_data = 0;
12'd4039: rgb_data = 0;
12'd4040: rgb_data = 0;
12'd4041: rgb_data = 0;
12'd4042: rgb_data = 0;
12'd4043: rgb_data = 0;
12'd4044: rgb_data = 0;
12'd4045: rgb_data = 0;
12'd4046: rgb_data = 0;
12'd4047: rgb_data = 0;
12'd4048: rgb_data = 0;
12'd4049: rgb_data = 0;
12'd4050: rgb_data = 0;
12'd4051: rgb_data = 0;
12'd4052: rgb_data = 0;
12'd4053: rgb_data = 0;
12'd4054: rgb_data = 0;
12'd4055: rgb_data = 0;
12'd4056: rgb_data = 0;
12'd4057: rgb_data = 0;
12'd4058: rgb_data = 0;
12'd4059: rgb_data = 0;
12'd4060: rgb_data = 0;
12'd4061: rgb_data = 0;
12'd4062: rgb_data = 0;
12'd4063: rgb_data = 0;
12'd4064: rgb_data = 0;
12'd4065: rgb_data = 0;
12'd4066: rgb_data = 0;
12'd4067: rgb_data = 0;
12'd4068: rgb_data = 0;
12'd4069: rgb_data = 0;
12'd4070: rgb_data = 0;
12'd4071: rgb_data = 0;
12'd4072: rgb_data = 0;
12'd4073: rgb_data = 0;
12'd4074: rgb_data = 0;
12'd4075: rgb_data = 0;
12'd4076: rgb_data = 0;
12'd4077: rgb_data = 0;
12'd4078: rgb_data = 0;
12'd4079: rgb_data = 0;
12'd4080: rgb_data = 0;
12'd4081: rgb_data = 0;
12'd4082: rgb_data = 0;
12'd4083: rgb_data = 0;
12'd4084: rgb_data = 0;
12'd4085: rgb_data = 0;
12'd4086: rgb_data = 0;
12'd4087: rgb_data = 0;
12'd4088: rgb_data = 0;
12'd4089: rgb_data = 0;
12'd4090: rgb_data = 0;
12'd4091: rgb_data = 0;
12'd4092: rgb_data = 0;
12'd4093: rgb_data = 0;
12'd4094: rgb_data = 0;
12'd4095: rgb_data = 0;

default : rgb_data = 8'd0;
endcase
endmodule
